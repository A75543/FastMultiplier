magic
tech scmos
timestamp 1715207069
<< polycontact >>
rect 115 270 119 274
rect 131 270 135 274
rect 147 270 151 274
rect 163 270 167 274
rect 179 270 183 274
rect 195 270 199 274
rect 211 270 215 274
rect 227 270 231 274
rect 2 20 6 24
rect -1106 -6 -1102 -2
rect -1090 -6 -1086 -2
rect -1074 -6 -1070 -2
rect -1058 -6 -1054 -2
rect -1042 -6 -1038 -2
rect -1026 -6 -1022 -2
rect -1010 -6 -1006 -2
rect -994 -6 -990 -2
<< metal1 >>
rect 113 302 115 306
rect 113 246 115 250
rect -4 56 0 60
rect -1219 40 -972 44
rect -968 24 2 28
rect -12 0 0 4
rect 14 -16 34 -12
rect 247 -84 282 -80
rect 6 -92 1195 -88
rect 46 -100 1059 -96
rect 86 -108 923 -104
rect 126 -116 787 -112
rect 166 -124 651 -120
rect 206 -132 515 -128
rect 246 -140 379 -136
rect -20 -220 -8 -216
rect -12 -276 0 -272
rect -22 -300 22 -296
rect -1183 -368 -16 -364
rect -158 -420 26 -416
rect -294 -556 30 -552
rect -430 -692 30 -688
rect -566 -828 30 -824
rect -702 -964 30 -960
rect -838 -1100 30 -1096
rect -974 -1236 30 -1232
rect 280 -2849 292 -2845
rect 288 -2913 292 -2909
rect 304 -2977 526 -2973
rect 312 -2985 810 -2981
rect 320 -2993 1322 -2989
rect 328 -3001 1834 -2997
rect 336 -3009 2346 -3005
rect 344 -3017 2858 -3013
rect 352 -3025 3370 -3021
rect 360 -3033 3882 -3029
rect 368 -3041 4162 -3037
rect 376 -3049 4442 -3045
rect 384 -3057 4722 -3053
rect 392 -3065 5002 -3061
rect 400 -3073 5282 -3069
rect 408 -3081 5442 -3077
rect 532 -3089 5466 -3085
rect 280 -3161 518 -3157
rect 288 -3217 526 -3213
rect 14 -3353 374 -3349
rect -12 -3361 358 -3357
<< m2contact >>
rect -8 56 -4 60
rect -1223 40 -1219 44
rect -972 40 -968 44
rect -972 24 -968 28
rect 2 24 6 28
rect -16 0 -12 4
rect 10 -16 14 -12
rect 243 -84 247 -80
rect 282 -84 286 -80
rect 2 -92 6 -88
rect 1195 -92 1199 -88
rect 42 -100 46 -96
rect 1059 -100 1063 -96
rect 82 -108 86 -104
rect 923 -108 927 -104
rect 122 -116 126 -112
rect 787 -116 791 -112
rect 162 -124 166 -120
rect 651 -124 655 -120
rect 202 -132 206 -128
rect 515 -132 519 -128
rect 242 -140 246 -136
rect 379 -140 383 -136
rect -1223 -256 -1219 -252
rect -26 -300 -22 -296
rect 22 -300 26 -296
rect -1187 -368 -1183 -364
rect -16 -368 -12 -364
rect -162 -420 -158 -416
rect -298 -556 -294 -552
rect -434 -692 -430 -688
rect -570 -828 -566 -824
rect -706 -964 -702 -960
rect -842 -1100 -838 -1096
rect -978 -1236 -974 -1232
rect 276 -2849 280 -2845
rect 526 -2889 530 -2885
rect 810 -2889 814 -2885
rect 1322 -2889 1326 -2885
rect 1834 -2889 1838 -2885
rect 2346 -2889 2350 -2885
rect 2858 -2889 2862 -2885
rect 3370 -2889 3374 -2885
rect 3882 -2889 3886 -2885
rect 4162 -2889 4166 -2885
rect 4442 -2889 4446 -2885
rect 4722 -2889 4726 -2885
rect 5002 -2889 5006 -2885
rect 5282 -2889 5286 -2885
rect 5442 -2889 5446 -2885
rect 284 -2913 288 -2909
rect 292 -2969 296 -2965
rect 300 -2977 304 -2973
rect 526 -2977 530 -2973
rect 308 -2985 312 -2981
rect 810 -2985 814 -2981
rect 316 -2993 320 -2989
rect 1322 -2993 1326 -2989
rect 324 -3001 328 -2997
rect 1834 -3001 1838 -2997
rect 332 -3009 336 -3005
rect 2346 -3009 2350 -3005
rect 5466 -3012 5470 -3008
rect 340 -3017 344 -3013
rect 2858 -3017 2862 -3013
rect 348 -3025 352 -3021
rect 3370 -3025 3374 -3021
rect 356 -3033 360 -3029
rect 3882 -3033 3886 -3029
rect 364 -3041 368 -3037
rect 4162 -3041 4166 -3037
rect 372 -3049 376 -3045
rect 4442 -3049 4446 -3045
rect 380 -3057 384 -3053
rect 4722 -3057 4726 -3053
rect 388 -3065 392 -3061
rect 5002 -3065 5006 -3061
rect 396 -3073 400 -3069
rect 5282 -3073 5286 -3069
rect 404 -3081 408 -3077
rect 5442 -3081 5446 -3077
rect 528 -3089 532 -3085
rect 5466 -3089 5470 -3085
rect 276 -3161 280 -3157
rect 284 -3217 288 -3213
rect 430 -3329 434 -3325
rect 10 -3353 14 -3349
rect -16 -3361 -12 -3357
rect 656 -3451 660 -3447
rect 792 -3451 796 -3447
rect 928 -3451 932 -3447
rect 1064 -3451 1068 -3447
rect 1200 -3451 1204 -3447
rect 1336 -3451 1340 -3447
rect 1472 -3451 1476 -3447
rect 1608 -3451 1612 -3447
rect 656 -3903 660 -3899
rect 792 -3903 796 -3899
rect 928 -3903 932 -3899
rect 1064 -3903 1068 -3899
rect 1200 -3903 1204 -3899
rect 1336 -3903 1340 -3899
rect 1472 -3903 1476 -3899
rect 1608 -3903 1612 -3899
<< metal2 >>
rect -1223 -252 -1219 40
rect -972 28 -968 40
rect -16 -276 -12 0
rect -8 -216 -4 56
rect 2 -248 6 -92
rect -1187 -364 -1183 -292
rect -978 -1232 -974 -300
rect -842 -1096 -838 -300
rect -706 -960 -702 -300
rect -570 -824 -566 -300
rect -434 -688 -430 -300
rect -298 -552 -294 -300
rect -162 -416 -158 -296
rect -16 -3357 -12 -368
rect 10 -3349 14 -16
rect 243 -80 247 -24
rect 42 -248 46 -100
rect 82 -248 86 -108
rect 122 -248 126 -116
rect 162 -248 166 -124
rect 202 -248 206 -132
rect 242 -248 246 -140
rect 282 -248 286 -84
rect 379 -136 383 -24
rect 515 -128 519 -24
rect 651 -120 655 -24
rect 787 -112 791 -24
rect 923 -104 927 -16
rect 1059 -96 1063 -8
rect 1195 -88 1199 -24
rect 22 -296 26 -280
rect 276 -3157 280 -2849
rect 284 -3213 288 -2913
rect 292 -3089 296 -2969
rect 526 -2973 530 -2889
rect 300 -3089 304 -2977
rect 810 -2981 814 -2889
rect 308 -3089 312 -2985
rect 1322 -2989 1326 -2889
rect 316 -3089 320 -2993
rect 1834 -2997 1838 -2889
rect 324 -3089 328 -3001
rect 2346 -3005 2350 -2889
rect 332 -3089 336 -3009
rect 2858 -3013 2862 -2889
rect 340 -3089 344 -3017
rect 3370 -3021 3374 -2889
rect 348 -3089 352 -3025
rect 3882 -3029 3886 -2889
rect 356 -3089 360 -3033
rect 364 -3089 368 -3041
rect 372 -3089 376 -3049
rect 4722 -3053 4726 -3040
rect 380 -3089 384 -3057
rect 5002 -3061 5006 -3032
rect 388 -3089 392 -3065
rect 5282 -3069 5286 -3024
rect 396 -3089 400 -3073
rect 5442 -3077 5446 -3016
rect 404 -3089 408 -3081
rect 5466 -3085 5470 -3012
rect 528 -3145 532 -3097
rect 544 -3145 548 -3141
rect 560 -3145 564 -3141
rect 576 -3145 580 -3141
rect 592 -3145 596 -3141
rect 608 -3145 612 -3141
rect 624 -3145 628 -3141
<< metal3 >>
rect -1220 312 5472 318
rect -1220 -4008 276 -4002
rect 287 -4008 5472 -4002
use 2Comp  2Comp_0
timestamp 1714367186
transform 1 0 113 0 1 246
box -117 -330 1096 66
use 2Comp  2Comp_1
timestamp 1714367186
transform 1 0 -1108 0 1 -30
box -117 -330 1096 66
use 16Bit2Complement  16Bit2Complement_0
timestamp 1714422570
transform 1 0 526 0 1 -3463
box -234 -536 1096 374
use MULT  MULT_0
timestamp 1714372070
transform 1 0 0 0 1 -1228
box -8 -1828 5472 1076
<< labels >>
rlabel metal1 114 248 114 248 1 VSS
rlabel polycontact 4 22 4 22 1 Sign
rlabel polycontact 117 272 117 272 1 A0
rlabel polycontact 133 272 133 272 1 A1
rlabel polycontact 149 272 149 272 1 A2
rlabel polycontact 165 272 165 272 1 A3
rlabel polycontact 181 272 181 272 1 A4
rlabel polycontact 197 272 197 272 1 A5
rlabel polycontact 213 272 213 272 1 A6
rlabel polycontact 229 272 229 272 1 A7
rlabel polycontact -1104 -4 -1104 -4 1 B0
rlabel polycontact -1088 -4 -1088 -4 1 B1
rlabel polycontact -1072 -4 -1072 -4 1 B2
rlabel polycontact -1056 -4 -1056 -4 1 B3
rlabel polycontact -1040 -4 -1040 -4 1 B4
rlabel polycontact -1024 -4 -1024 -4 1 B5
rlabel polycontact -1008 -4 -1008 -4 1 B6
rlabel polycontact -992 -4 -992 -4 1 B7
rlabel metal1 114 304 114 304 1 VDD
rlabel m2contact 432 -3327 432 -3327 1 XOR
rlabel m2contact 1610 -3901 1610 -3901 1 Q15
rlabel m2contact 1474 -3901 1474 -3901 1 Q14
rlabel m2contact 1338 -3901 1338 -3901 1 Q13
rlabel m2contact 1202 -3901 1202 -3901 1 Q12
rlabel m2contact 1066 -3901 1066 -3901 1 Q11
rlabel m2contact 930 -3901 930 -3901 1 Q10
rlabel m2contact 794 -3901 794 -3901 1 Q9
rlabel m2contact 658 -3901 658 -3901 1 Q8
rlabel m2contact 1610 -3449 1610 -3449 1 Q7
rlabel m2contact 1474 -3449 1474 -3449 1 Q6
rlabel m2contact 1338 -3449 1338 -3449 1 Q5
rlabel m2contact 1202 -3449 1202 -3449 1 Q4
rlabel m2contact 1066 -3449 1066 -3449 1 Q3
rlabel m2contact 930 -3449 930 -3449 1 Q2
rlabel m2contact 794 -3449 794 -3449 1 Q1
rlabel m2contact 658 -3449 658 -3449 1 Q0
rlabel m2contact 5468 -3010 5468 -3010 1 q0
rlabel m2contact 5444 -2887 5444 -2887 1 q1
rlabel m2contact 5284 -2887 5284 -2887 1 q2
rlabel m2contact 5004 -2887 5004 -2887 1 q3
rlabel m2contact 4724 -2887 4724 -2887 1 q4
rlabel m2contact 4444 -2887 4444 -2887 1 q5
rlabel m2contact 4164 -2887 4164 -2887 1 q6
rlabel m2contact 3884 -2887 3884 -2887 1 q7
rlabel m2contact 3372 -2887 3372 -2887 1 q8
rlabel m2contact 2860 -2887 2860 -2887 1 q9
rlabel m2contact 2348 -2887 2348 -2887 1 q10
rlabel m2contact 1836 -2887 1836 -2887 1 q11
rlabel m2contact 1324 -2887 1324 -2887 1 q12
rlabel m2contact 812 -2887 812 -2887 1 q13
rlabel m2contact 528 -2887 528 -2887 1 q14
rlabel m2contact 294 -2967 294 -2967 1 q15
<< end >>
