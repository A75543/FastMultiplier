magic
tech scmos
timestamp 1714291806
<< polycontact >>
rect 18 -96 22 -92
<< metal1 >>
rect -4 56 0 60
rect -68 20 2 24
rect 128 0 1092 4
rect -12 -8 114 -4
rect 126 -8 841 -4
rect -20 -16 98 -12
rect 110 -16 721 -12
rect -28 -24 82 -20
rect 94 -24 601 -20
rect -36 -32 66 -28
rect 78 -32 481 -28
rect -44 -40 50 -36
rect 62 -40 361 -36
rect -52 -48 34 -44
rect 46 -48 242 -44
rect -60 -56 18 -52
rect 30 -56 122 -52
rect -4 -64 0 -60
rect 959 -128 1092 -124
rect 62 -176 114 -172
rect 198 -176 234 -172
rect 334 -176 354 -172
rect 470 -176 473 -172
rect 597 -176 602 -172
rect 717 -176 738 -172
rect 837 -176 874 -172
rect 957 -176 1010 -172
rect -4 -190 0 -186
rect 1088 -246 1092 -242
rect 6 -262 10 -258
rect -12 -274 970 -270
rect -20 -282 834 -278
rect -28 -290 698 -286
rect -36 -298 562 -294
rect -44 -306 426 -302
rect -52 -314 290 -310
rect -60 -322 154 -318
rect -68 -330 18 -326
<< m2contact >>
rect -8 56 -4 60
rect -72 20 -68 24
rect 2 20 6 24
rect 18 20 22 24
rect 34 20 38 24
rect 50 20 54 24
rect 66 20 70 24
rect 82 20 86 24
rect 98 20 102 24
rect 114 20 118 24
rect 10 12 14 16
rect 26 12 30 16
rect 42 12 46 16
rect 58 12 62 16
rect 74 12 78 16
rect 90 12 94 16
rect 106 12 110 16
rect 122 12 126 16
rect 1092 0 1096 4
rect -16 -8 -12 -4
rect 114 -8 118 -4
rect 122 -8 126 -4
rect 841 -8 845 -4
rect -24 -16 -20 -12
rect 98 -16 102 -12
rect 106 -16 110 -12
rect 721 -16 725 -12
rect -32 -24 -28 -20
rect 82 -24 86 -20
rect 90 -24 94 -20
rect 601 -24 605 -20
rect -40 -32 -36 -28
rect 66 -32 70 -28
rect 74 -32 78 -28
rect 481 -32 485 -28
rect -48 -40 -44 -36
rect 50 -40 54 -36
rect 58 -40 62 -36
rect 361 -40 365 -36
rect -56 -48 -52 -44
rect 34 -48 38 -44
rect 42 -48 46 -44
rect 242 -48 246 -44
rect -64 -56 -60 -52
rect 18 -56 22 -52
rect 26 -56 30 -52
rect 122 -56 126 -52
rect -8 -64 -4 -60
rect 122 -92 126 -88
rect 242 -92 246 -88
rect 361 -92 365 -88
rect 481 -92 485 -88
rect 601 -92 605 -88
rect 721 -92 725 -88
rect 841 -92 845 -88
rect 114 -108 118 -104
rect 234 -108 238 -104
rect 354 -108 358 -104
rect 473 -108 477 -104
rect 593 -108 597 -104
rect 713 -108 717 -104
rect 833 -108 837 -104
rect 953 -108 957 -104
rect 1092 -128 1096 -124
rect 10 -144 14 -140
rect 58 -176 62 -172
rect 114 -176 118 -172
rect 194 -176 198 -172
rect 234 -176 238 -172
rect 330 -176 334 -172
rect 354 -176 358 -172
rect 466 -176 470 -172
rect 473 -176 477 -172
rect 593 -176 597 -172
rect 602 -176 606 -172
rect 713 -176 717 -172
rect 738 -176 742 -172
rect 833 -176 837 -172
rect 874 -176 878 -172
rect 953 -176 957 -172
rect 1010 -176 1014 -172
rect -8 -190 -4 -186
rect 130 -234 134 -230
rect 266 -234 270 -230
rect 402 -234 406 -230
rect 538 -234 542 -230
rect 674 -234 678 -230
rect 810 -234 814 -230
rect 946 -234 950 -230
rect 1082 -234 1086 -230
rect 1092 -246 1096 -242
rect -16 -274 -12 -270
rect 970 -274 974 -270
rect -24 -282 -20 -278
rect 834 -282 838 -278
rect -32 -290 -28 -286
rect 698 -290 702 -286
rect -40 -298 -36 -294
rect 562 -298 566 -294
rect -48 -306 -44 -302
rect 426 -306 430 -302
rect -56 -314 -52 -310
rect 290 -314 294 -310
rect -64 -322 -60 -318
rect 154 -322 158 -318
rect -72 -330 -68 -326
rect 18 -330 22 -326
<< metal2 >>
rect -72 -326 -68 20
rect -64 -318 -60 -56
rect -56 -310 -52 -48
rect -48 -302 -44 -40
rect -40 -294 -36 -32
rect -32 -286 -28 -24
rect -24 -278 -20 -16
rect -16 -270 -12 -8
rect -8 -60 -4 56
rect -8 -186 -4 -64
rect 10 -140 14 12
rect 18 -52 22 20
rect 26 -52 30 12
rect 34 -44 38 20
rect 42 -44 46 12
rect 50 -36 54 20
rect 58 -36 62 12
rect 66 -28 70 20
rect 74 -28 78 12
rect 82 -20 86 20
rect 90 -20 94 12
rect 98 -12 102 20
rect 106 -12 110 12
rect 114 -4 118 20
rect 122 -4 126 12
rect 122 -88 126 -56
rect 242 -88 246 -48
rect 361 -88 365 -40
rect 481 -88 485 -32
rect 601 -88 605 -24
rect 721 -88 725 -16
rect 841 -88 845 -8
rect 18 -96 22 -92
rect 114 -172 118 -108
rect 234 -172 238 -108
rect 354 -172 358 -108
rect 473 -172 477 -108
rect 593 -172 597 -108
rect 713 -172 717 -108
rect 833 -172 837 -108
rect 953 -172 957 -108
rect 1092 -124 1096 0
rect 58 -218 62 -176
rect 194 -218 198 -176
rect 330 -218 334 -176
rect 466 -218 470 -176
rect 602 -218 606 -176
rect 738 -218 742 -176
rect 874 -218 878 -176
rect 1010 -218 1014 -176
rect 1092 -242 1096 -128
rect 18 -326 22 -270
rect 154 -318 158 -270
rect 290 -310 294 -270
rect 426 -302 430 -270
rect 562 -294 566 -270
rect 698 -286 702 -270
rect 834 -278 838 -270
use 8bitAdder  8bitAdder_0
timestamp 1714184300
transform 1 0 0 0 1 -128
box -4 -40 961 71
use 8bitINV  8bitINV_0
timestamp 1711614163
transform 1 0 0 0 1 0
box -4 0 132 66
use mux2x1_8  mux2x1_8_0
timestamp 1711616816
transform 1 0 0 0 1 -246
box -4 -24 1094 66
<< labels >>
rlabel metal2 20 -94 20 -94 1 B
rlabel metal1 8 -260 8 -260 1 S
rlabel m2contact 132 -232 132 -232 1 Y0
rlabel m2contact 268 -232 268 -232 1 Y1
rlabel m2contact 404 -232 404 -232 1 Y2
rlabel m2contact 540 -232 540 -232 1 Y3
rlabel m2contact 676 -232 676 -232 1 Y4
rlabel m2contact 812 -232 812 -232 1 Y5
rlabel m2contact 948 -232 948 -232 1 Y6
rlabel m2contact 1084 -232 1084 -232 1 Y7
rlabel metal1 -2 58 -2 58 1 VDD
rlabel metal1 130 2 130 2 1 VSS
rlabel m2contact 4 22 4 22 1 A0
rlabel m2contact 20 22 20 22 1 A1
rlabel m2contact 36 22 36 22 1 A2
rlabel m2contact 52 22 52 22 1 A3
rlabel m2contact 68 22 68 22 1 A4
rlabel m2contact 84 22 84 22 1 A5
rlabel m2contact 100 22 100 22 1 A6
rlabel m2contact 116 22 116 22 1 A7
<< end >>
