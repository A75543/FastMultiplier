magic
tech scmos
timestamp 1711067998
<< nwell >>
rect -36 38 50 71
<< ntransistor >>
rect -25 8 -23 12
rect -9 8 -7 12
rect 7 8 9 12
rect 15 8 17 12
rect 23 8 25 12
rect 31 8 33 12
<< ptransistor >>
rect -25 44 -23 52
rect -9 44 -7 52
rect 7 44 9 52
rect 15 44 17 52
rect 23 44 25 52
rect 31 44 33 52
<< ndiffusion >>
rect -26 8 -25 12
rect -23 8 -22 12
rect -10 8 -9 12
rect -7 8 -6 12
rect 6 8 7 12
rect 9 8 15 12
rect 17 8 18 12
rect 22 8 23 12
rect 25 8 31 12
rect 33 8 34 12
<< pdiffusion >>
rect -26 44 -25 52
rect -23 44 -22 52
rect -10 44 -9 52
rect -7 44 -6 52
rect 6 44 7 52
rect 9 44 10 52
rect 14 44 15 52
rect 17 44 18 52
rect 22 44 23 52
rect 25 44 26 52
rect 30 44 31 52
rect 33 44 34 52
<< ndcontact >>
rect -30 8 -26 12
rect -22 8 -18 12
rect -14 8 -10 12
rect -6 8 -2 12
rect 2 8 6 12
rect 18 8 22 12
rect 34 8 38 12
<< pdcontact >>
rect -30 44 -26 52
rect -22 44 -18 52
rect -14 44 -10 52
rect -6 44 -2 52
rect 2 44 6 52
rect 10 44 14 52
rect 18 44 22 52
rect 26 44 30 52
rect 34 44 38 52
<< psubstratepcontact >>
rect -30 0 -26 4
rect -14 0 -10 4
rect 18 0 22 4
<< nsubstratencontact >>
rect -30 64 -26 68
rect -14 64 -10 68
rect 10 64 14 68
<< polysilicon >>
rect -25 52 -23 54
rect -9 52 -7 54
rect 7 52 9 54
rect 15 52 17 54
rect 23 52 25 54
rect 31 52 33 54
rect -25 28 -23 44
rect -9 28 -7 44
rect 7 28 9 44
rect 15 28 17 44
rect 23 32 25 44
rect -26 24 -23 28
rect -10 24 -7 28
rect 6 24 9 28
rect 16 24 17 28
rect 20 28 25 32
rect 24 24 25 28
rect -25 12 -23 24
rect -9 12 -7 24
rect 7 12 9 24
rect 15 12 17 24
rect 23 12 25 24
rect 31 32 33 44
rect 31 28 35 32
rect 31 12 33 24
rect -25 6 -23 8
rect -9 6 -7 8
rect 7 6 9 8
rect 15 6 17 8
rect 23 6 25 8
rect 31 6 33 8
<< polycontact >>
rect -30 24 -26 28
rect -14 24 -10 28
rect 2 24 6 28
rect 12 24 16 28
rect 20 24 24 28
rect 31 24 35 28
<< metal1 >>
rect -32 64 -30 68
rect -26 64 -14 68
rect -10 64 10 68
rect 14 64 48 68
rect -30 52 -26 64
rect -14 52 -10 64
rect 10 52 14 64
rect -22 16 -18 44
rect -6 16 -2 44
rect 18 56 38 60
rect 18 52 22 56
rect 34 52 38 56
rect 2 40 6 44
rect 18 40 22 44
rect 2 36 22 40
rect 26 40 30 44
rect 26 36 46 40
rect 42 20 46 36
rect 2 16 46 20
rect 2 12 6 16
rect 34 12 38 16
rect -30 4 -26 8
rect -14 4 -10 8
rect 18 4 22 8
rect -32 0 -30 4
rect -26 0 -14 4
rect -10 0 18 4
rect 22 0 48 4
rect -10 -8 12 -4
rect -26 -16 2 -12
rect -18 -24 20 -20
rect -2 -32 31 -28
<< m2contact >>
rect -30 28 -26 32
rect -14 28 -10 32
rect -22 12 -18 16
rect 2 28 6 32
rect 12 28 16 32
rect 20 28 24 32
rect 31 28 35 32
rect -6 12 -2 16
rect -14 -8 -10 -4
rect 12 -8 16 -4
rect -30 -16 -26 -12
rect 2 -16 6 -12
rect -22 -24 -18 -20
rect 20 -24 24 -20
rect -6 -32 -2 -28
rect 31 -32 35 -28
<< metal2 >>
rect -30 -12 -26 28
rect -22 -20 -18 12
rect -14 -4 -10 28
rect -6 -28 -2 12
rect 2 -12 6 28
rect 12 -4 16 28
rect 20 -20 24 28
rect 31 -28 35 28
<< labels >>
rlabel psubstratepcontact 20 2 20 2 1 VSS
rlabel psubstratepcontact -12 2 -12 2 1 VSS
rlabel psubstratepcontact -28 2 -28 2 1 VSS
rlabel metal1 44 26 44 26 1 Y
rlabel nsubstratencontact 12 66 12 66 1 VDD
rlabel nsubstratencontact -28 66 -28 66 1 VDD
rlabel nsubstratencontact -12 66 -12 66 1 VDD
rlabel polycontact -12 26 -12 26 1 B
rlabel polycontact -28 26 -28 26 1 A
<< end >>
