magic
tech scmos
timestamp 1714342102
<< metal1 >>
rect -4 56 0 60
rect 320 0 324 4
rect 26 -8 30 -4
rect -4 -80 0 -76
rect 320 -136 324 -132
rect 26 -144 30 -140
rect -4 -216 0 -212
rect 320 -272 324 -268
rect 26 -280 30 -276
rect -4 -352 0 -348
rect 320 -408 324 -404
rect 26 -416 30 -412
rect -4 -488 0 -484
rect 320 -544 324 -540
rect 26 -552 30 -548
rect -4 -624 0 -620
rect 320 -680 324 -676
rect 26 -688 30 -684
rect -4 -760 0 -756
rect 320 -816 324 -812
rect 26 -824 30 -820
rect -4 -896 0 -892
rect 320 -952 324 -948
rect 26 -960 30 -956
<< m2contact >>
rect 34 120 38 124
rect 74 112 78 116
rect 114 104 118 108
rect 154 96 158 100
rect 194 88 198 92
rect 234 80 238 84
rect 274 72 278 76
rect 314 64 318 68
rect -8 56 -4 60
rect 2 24 6 28
rect 42 24 46 28
rect 82 24 86 28
rect 122 24 126 28
rect 162 24 166 28
rect 202 24 206 28
rect 242 24 246 28
rect 282 24 286 28
rect 324 0 328 4
rect 34 -16 38 -12
rect 74 -24 78 -20
rect 114 -32 118 -28
rect 154 -40 158 -36
rect 194 -48 198 -44
rect 234 -56 238 -52
rect 274 -64 278 -60
rect 314 -72 318 -68
rect -8 -80 -4 -76
rect 2 -112 6 -108
rect 42 -112 46 -108
rect 82 -112 86 -108
rect 122 -112 126 -108
rect 162 -112 166 -108
rect 202 -112 206 -108
rect 242 -112 246 -108
rect 282 -112 286 -108
rect 324 -136 328 -132
rect 34 -152 38 -148
rect 74 -160 78 -156
rect 114 -168 118 -164
rect 154 -176 158 -172
rect 194 -184 198 -180
rect 234 -192 238 -188
rect 274 -200 278 -196
rect 314 -208 318 -204
rect -8 -216 -4 -212
rect 2 -248 6 -244
rect 42 -248 46 -244
rect 82 -248 86 -244
rect 122 -248 126 -244
rect 162 -248 166 -244
rect 202 -248 206 -244
rect 242 -248 246 -244
rect 282 -248 286 -244
rect 324 -272 328 -268
rect 34 -288 38 -284
rect 74 -296 78 -292
rect 114 -304 118 -300
rect 154 -312 158 -308
rect 194 -320 198 -316
rect 234 -328 238 -324
rect 274 -336 278 -332
rect 314 -344 318 -340
rect -8 -352 -4 -348
rect 2 -384 6 -380
rect 42 -384 46 -380
rect 82 -384 86 -380
rect 122 -384 126 -380
rect 162 -384 166 -380
rect 202 -384 206 -380
rect 242 -384 246 -380
rect 282 -384 286 -380
rect 324 -408 328 -404
rect 34 -424 38 -420
rect 74 -432 78 -428
rect 114 -440 118 -436
rect 154 -448 158 -444
rect 194 -456 198 -452
rect 234 -464 238 -460
rect 274 -472 278 -468
rect 314 -480 318 -476
rect -8 -488 -4 -484
rect 2 -520 6 -516
rect 42 -520 46 -516
rect 82 -520 86 -516
rect 122 -520 126 -516
rect 162 -520 166 -516
rect 202 -520 206 -516
rect 242 -520 246 -516
rect 282 -520 286 -516
rect 324 -544 328 -540
rect 34 -560 38 -556
rect 74 -568 78 -564
rect 114 -576 118 -572
rect 154 -584 158 -580
rect 194 -592 198 -588
rect 234 -600 238 -596
rect 274 -608 278 -604
rect 314 -616 318 -612
rect -8 -624 -4 -620
rect 2 -656 6 -652
rect 42 -656 46 -652
rect 82 -656 86 -652
rect 122 -656 126 -652
rect 162 -656 166 -652
rect 202 -656 206 -652
rect 242 -656 246 -652
rect 282 -656 286 -652
rect 324 -680 328 -676
rect 34 -696 38 -692
rect 74 -704 78 -700
rect 114 -712 118 -708
rect 154 -720 158 -716
rect 194 -728 198 -724
rect 234 -736 238 -732
rect 274 -744 278 -740
rect 314 -752 318 -748
rect -8 -760 -4 -756
rect 2 -792 6 -788
rect 42 -792 46 -788
rect 82 -792 86 -788
rect 122 -792 126 -788
rect 162 -792 166 -788
rect 202 -792 206 -788
rect 242 -792 246 -788
rect 282 -792 286 -788
rect 324 -816 328 -812
rect 34 -832 38 -828
rect 74 -840 78 -836
rect 114 -848 118 -844
rect 154 -856 158 -852
rect 194 -864 198 -860
rect 234 -872 238 -868
rect 274 -880 278 -876
rect 314 -888 318 -884
rect -8 -896 -4 -892
rect 2 -928 6 -924
rect 42 -928 46 -924
rect 82 -928 86 -924
rect 122 -928 126 -924
rect 162 -928 166 -924
rect 202 -928 206 -924
rect 242 -928 246 -924
rect 282 -928 286 -924
rect 324 -952 328 -948
<< metal2 >>
rect -8 -76 -4 56
rect -8 -212 -4 -80
rect -8 -348 -4 -216
rect -8 -484 -4 -352
rect -8 -620 -4 -488
rect -8 -756 -4 -624
rect -8 -892 -4 -760
rect 2 -108 6 24
rect 2 -244 6 -112
rect 42 -108 46 24
rect 2 -380 6 -248
rect 42 -244 46 -112
rect 82 -108 86 24
rect 2 -516 6 -384
rect 42 -380 46 -248
rect 82 -244 86 -112
rect 122 -108 126 24
rect 2 -652 6 -520
rect 42 -516 46 -384
rect 82 -380 86 -248
rect 122 -244 126 -112
rect 162 -108 166 24
rect 2 -788 6 -656
rect 42 -652 46 -520
rect 82 -516 86 -384
rect 122 -380 126 -248
rect 162 -244 166 -112
rect 202 -108 206 24
rect 2 -924 6 -792
rect 42 -788 46 -656
rect 82 -652 86 -520
rect 122 -516 126 -384
rect 162 -380 166 -248
rect 202 -244 206 -112
rect 242 -108 246 24
rect 42 -924 46 -792
rect 82 -788 86 -656
rect 122 -652 126 -520
rect 162 -516 166 -384
rect 202 -380 206 -248
rect 242 -244 246 -112
rect 282 -108 286 24
rect 82 -924 86 -792
rect 122 -788 126 -656
rect 162 -652 166 -520
rect 202 -516 206 -384
rect 242 -380 246 -248
rect 282 -244 286 -112
rect 324 -132 328 0
rect 122 -924 126 -792
rect 162 -788 166 -656
rect 202 -652 206 -520
rect 242 -516 246 -384
rect 282 -380 286 -248
rect 324 -268 328 -136
rect 162 -924 166 -792
rect 202 -788 206 -656
rect 242 -652 246 -520
rect 282 -516 286 -384
rect 324 -404 328 -272
rect 202 -924 206 -792
rect 242 -788 246 -656
rect 282 -652 286 -520
rect 324 -540 328 -408
rect 242 -924 246 -792
rect 282 -788 286 -656
rect 324 -676 328 -544
rect 282 -924 286 -792
rect 324 -812 328 -680
rect 324 -948 328 -816
use 8bitAND  8bitAND_0
timestamp 1714340751
transform 1 0 0 0 1 0
box -4 -8 892 124
use 8bitAND  8bitAND_1
timestamp 1714340751
transform 1 0 0 0 1 -136
box -4 -8 892 124
use 8bitAND  8bitAND_2
timestamp 1714340751
transform 1 0 0 0 1 -272
box -4 -8 892 124
use 8bitAND  8bitAND_3
timestamp 1714340751
transform 1 0 0 0 1 -408
box -4 -8 892 124
use 8bitAND  8bitAND_4
timestamp 1714340751
transform 1 0 0 0 1 -544
box -4 -8 892 124
use 8bitAND  8bitAND_5
timestamp 1714340751
transform 1 0 0 0 1 -680
box -4 -8 892 124
use 8bitAND  8bitAND_6
timestamp 1714340751
transform 1 0 0 0 1 -816
box -4 -8 892 124
use 8bitAND  8bitAND_7
timestamp 1714340751
transform 1 0 0 0 1 -952
box -4 -8 892 124
<< labels >>
rlabel metal1 28 -6 28 -6 1 M7
rlabel m2contact 4 26 4 26 1 A7
rlabel m2contact 44 26 44 26 1 A6
rlabel m2contact 84 26 84 26 1 A5
rlabel m2contact 124 26 124 26 1 A4
rlabel m2contact 164 26 164 26 1 A3
rlabel m2contact 204 26 204 26 1 A2
rlabel m2contact 244 26 244 26 1 A1
rlabel m2contact 284 26 284 26 1 A0
rlabel metal1 322 2 322 2 1 VSS
rlabel metal1 28 -142 28 -142 1 M6
rlabel metal1 28 -278 28 -278 1 M5
rlabel metal1 28 -686 28 -686 1 M2
rlabel metal1 28 -822 28 -822 1 M1
rlabel metal1 28 -958 28 -958 1 M0
rlabel metal1 28 -414 28 -414 1 M4
rlabel metal1 28 -550 28 -550 1 M3
rlabel m2contact 36 122 36 122 5 P7_7
rlabel m2contact 76 114 76 114 1 P7_6
rlabel m2contact 116 106 116 106 1 P7_5
rlabel m2contact 156 98 156 98 1 P7_4
rlabel m2contact 196 90 196 90 1 P7_3
rlabel m2contact 236 82 236 82 1 P7_2
rlabel m2contact 276 74 276 74 1 P7_1
rlabel m2contact 316 66 316 66 1 P7_0
rlabel m2contact 36 -14 36 -14 1 P6_7
rlabel m2contact 76 -22 76 -22 1 P6_6
rlabel m2contact 116 -30 116 -30 1 P6_5
rlabel m2contact 156 -38 156 -38 1 P6_4
rlabel m2contact 196 -46 196 -46 1 P6_3
rlabel m2contact 236 -54 236 -54 1 P6_2
rlabel m2contact 276 -62 276 -62 1 P6_1
rlabel m2contact 316 -70 316 -70 1 P6_0
rlabel m2contact 36 -150 36 -150 1 P5_7
rlabel m2contact 76 -158 76 -158 1 P5_6
rlabel m2contact 116 -166 116 -166 1 P5_5
rlabel m2contact 156 -174 156 -174 1 P5_4
rlabel m2contact 196 -182 196 -182 1 P5_3
rlabel m2contact 236 -190 236 -190 1 P5_2
rlabel m2contact 276 -198 276 -198 1 P5_1
rlabel m2contact 316 -206 316 -206 1 P5_0
rlabel m2contact 36 -286 36 -286 1 P4_7
rlabel m2contact 76 -294 76 -294 1 P4_6
rlabel m2contact 116 -302 116 -302 1 P4_5
rlabel m2contact 156 -310 156 -310 1 P4_4
rlabel m2contact 196 -318 196 -318 1 P4_3
rlabel m2contact 236 -326 236 -326 1 P4_2
rlabel m2contact 276 -334 276 -334 1 P4_1
rlabel m2contact 316 -342 316 -342 1 P4_0
rlabel m2contact 36 -422 36 -422 1 P3_7
rlabel m2contact 76 -430 76 -430 1 P3_6
rlabel m2contact 116 -438 116 -438 1 P3_5
rlabel m2contact 157 -446 157 -446 1 P3_4
rlabel m2contact 196 -454 196 -454 1 P3_3
rlabel m2contact 236 -462 236 -462 1 P3_2
rlabel m2contact 276 -470 276 -470 1 P3_1
rlabel m2contact 316 -478 316 -478 1 P3_0
rlabel m2contact 36 -558 36 -558 1 P2_7
rlabel m2contact 76 -566 76 -566 1 P2_6
rlabel m2contact 116 -574 116 -574 1 P2_5
rlabel m2contact 156 -582 156 -582 1 P2_4
rlabel m2contact 196 -590 196 -590 1 P2_3
rlabel m2contact 236 -598 236 -598 1 P2_2
rlabel m2contact 276 -606 276 -606 1 P2_1
rlabel m2contact 316 -614 316 -614 1 P2_0
rlabel m2contact 36 -694 36 -694 1 P1_7
rlabel m2contact 76 -702 76 -702 1 P1_6
rlabel m2contact 116 -710 116 -710 1 P1_5
rlabel m2contact 156 -718 156 -718 1 P1_4
rlabel m2contact 196 -726 196 -726 1 P1_3
rlabel m2contact 236 -734 236 -734 1 P1_2
rlabel m2contact 276 -742 276 -742 1 P1_1
rlabel m2contact 316 -750 316 -750 1 P1_0
rlabel m2contact 36 -830 36 -830 1 P0_7
rlabel m2contact 76 -838 76 -838 1 P0_6
rlabel m2contact 116 -846 116 -846 1 P0_5
rlabel m2contact 156 -854 156 -854 1 P0_4
rlabel m2contact 196 -862 196 -862 1 P0_3
rlabel m2contact 236 -870 236 -870 1 P0_2
rlabel m2contact 276 -878 276 -878 1 P0_1
rlabel m2contact 316 -886 316 -886 1 P0_0
rlabel metal1 -2 58 -2 58 1 VDD
<< end >>
