magic
tech scmos
timestamp 1711614163
<< nwell >>
rect 0 56 2 60
<< polycontact >>
rect 2 24 6 28
rect 18 24 22 28
rect 34 24 38 28
rect 50 24 54 28
rect 66 24 70 28
rect 82 24 86 28
rect 98 24 102 28
rect 114 24 118 28
<< metal1 >>
rect 0 56 2 60
rect 10 24 14 28
rect 26 24 30 28
rect 42 24 46 28
rect 58 24 62 28
rect 74 24 78 28
rect 90 24 94 28
rect 106 24 110 28
rect 122 24 126 28
rect 0 0 2 4
use INV  INV_0
timestamp 1711614163
transform 1 0 0 0 1 0
box -4 0 20 66
use INV  INV_1
timestamp 1711614163
transform 1 0 16 0 1 0
box -4 0 20 66
use INV  INV_2
timestamp 1711614163
transform 1 0 32 0 1 0
box -4 0 20 66
use INV  INV_3
timestamp 1711614163
transform 1 0 48 0 1 0
box -4 0 20 66
use INV  INV_4
timestamp 1711614163
transform 1 0 64 0 1 0
box -4 0 20 66
use INV  INV_5
timestamp 1711614163
transform 1 0 80 0 1 0
box -4 0 20 66
use INV  INV_6
timestamp 1711614163
transform 1 0 96 0 1 0
box -4 0 20 66
use INV  INV_7
timestamp 1711614163
transform 1 0 112 0 1 0
box -4 0 20 66
<< labels >>
rlabel metal1 1 58 1 58 1 VDD
rlabel metal1 1 2 1 2 1 VSS
rlabel polycontact 4 26 4 26 1 A0
rlabel polycontact 20 26 20 26 1 A1
rlabel polycontact 36 26 36 26 1 A2
rlabel polycontact 52 26 52 26 1 A3
rlabel polycontact 68 26 68 26 1 A4
rlabel polycontact 84 26 84 26 1 A5
rlabel polycontact 100 26 100 26 1 A6
rlabel polycontact 116 26 116 26 1 A7
rlabel metal1 12 26 12 26 1 Y0
rlabel metal1 28 26 28 26 1 Y1
rlabel metal1 44 26 44 26 1 Y2
rlabel metal1 60 26 60 26 1 Y3
rlabel metal1 76 26 76 26 1 Y4
rlabel metal1 92 26 92 26 1 Y5
rlabel metal1 108 26 108 26 1 Y6
rlabel metal1 124 26 124 26 1 Y7
<< end >>
