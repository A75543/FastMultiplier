magic
tech scmos
timestamp 1711561704
<< nwell >>
rect -4 38 44 66
<< ntransistor >>
rect 7 8 9 16
rect 15 8 17 16
rect 31 8 33 16
<< ptransistor >>
rect 7 44 9 52
rect 15 44 17 52
rect 31 44 33 52
<< ndiffusion >>
rect 6 8 7 16
rect 9 8 15 16
rect 17 8 18 16
rect 30 8 31 16
rect 33 8 34 16
<< pdiffusion >>
rect 6 44 7 52
rect 9 44 10 52
rect 14 44 15 52
rect 17 44 18 52
rect 30 44 31 52
rect 33 44 34 52
<< ndcontact >>
rect 2 8 6 16
rect 18 8 22 16
rect 26 8 30 16
rect 34 8 38 16
<< pdcontact >>
rect 2 44 6 52
rect 10 44 14 52
rect 18 44 22 52
rect 26 44 30 52
rect 34 44 38 52
<< psubstratepcontact >>
rect 2 0 6 4
rect 26 0 30 4
<< nsubstratencontact >>
rect 2 56 6 60
rect 18 56 22 60
rect 26 56 30 60
<< polysilicon >>
rect 7 52 9 54
rect 15 52 17 54
rect 31 52 33 54
rect 7 24 9 44
rect 6 20 9 24
rect 7 16 9 20
rect 15 40 17 44
rect 15 36 18 40
rect 15 16 17 36
rect 31 16 33 44
rect 7 6 9 8
rect 15 6 17 8
rect 31 6 33 8
<< polycontact >>
rect 2 20 6 24
rect 18 36 22 40
rect 27 28 31 32
<< metal1 >>
rect 0 56 2 60
rect 6 56 18 60
rect 22 56 26 60
rect 30 56 40 60
rect 2 52 6 56
rect 18 52 22 56
rect 26 52 30 56
rect 10 32 14 44
rect 10 28 27 32
rect 18 16 22 28
rect 34 16 38 44
rect 2 4 6 8
rect 26 4 30 8
rect 0 0 2 4
rect 6 0 26 4
rect 30 0 40 4
<< labels >>
rlabel polycontact 4 22 4 22 3 A
rlabel psubstratepcontact 4 2 4 2 2 VSS
rlabel psubstratepcontact 28 2 28 2 1 VSS
rlabel nsubstratencontact 4 58 4 58 4 VDD
rlabel polycontact 20 38 20 38 7 B
rlabel nsubstratencontact 20 58 20 58 6 VDD
rlabel metal1 36 30 36 30 1 Y
rlabel nsubstratencontact 28 58 28 58 1 VDD
<< end >>
