magic
tech scmos
timestamp 1714372070
<< nwell >>
rect 343 -59 346 -55
<< metal1 >>
rect 849 1072 5472 1076
rect 849 1064 5472 1068
rect 849 1056 1870 1060
rect 1874 1056 5472 1060
rect 849 1048 2382 1052
rect 2386 1048 5472 1052
rect 849 1040 2894 1044
rect 2898 1040 5472 1044
rect 849 1032 3406 1036
rect 3410 1032 5472 1036
rect 849 1024 3918 1028
rect 3922 1024 5472 1028
rect 849 1016 5074 1020
rect 5078 1016 5472 1020
rect -4 1008 0 1012
rect 0 952 2 956
rect 26 944 30 948
rect 849 936 5472 940
rect 849 928 5472 932
rect 849 920 1878 924
rect 1882 920 5472 924
rect 849 912 2390 916
rect 2394 912 5472 916
rect 849 904 2902 908
rect 2906 904 5472 908
rect 849 896 3414 900
rect 3418 896 5472 900
rect 849 888 4430 892
rect 4434 888 5472 892
rect 849 880 4942 884
rect 4946 880 5472 884
rect 26 808 30 812
rect 849 800 5472 804
rect 849 792 922 796
rect 926 792 5472 796
rect 849 784 1886 788
rect 1890 784 5472 788
rect 849 776 2398 780
rect 2402 776 5472 780
rect 849 768 2910 772
rect 2914 768 5472 772
rect 849 760 3926 764
rect 3930 760 5472 764
rect 849 752 4438 756
rect 4442 752 5472 756
rect 849 744 4950 748
rect 4954 744 5472 748
rect 26 672 30 676
rect 849 664 906 668
rect 910 664 5472 668
rect 849 656 1202 660
rect 1206 656 5472 660
rect 849 648 1894 652
rect 1898 648 5472 652
rect 849 640 2406 644
rect 2410 640 5472 644
rect 849 632 3422 636
rect 3426 632 5472 636
rect 849 624 3934 628
rect 3938 624 5472 628
rect 849 616 4446 620
rect 4450 616 5472 620
rect 849 608 4958 612
rect 4962 608 5472 612
rect 26 536 30 540
rect 849 528 1186 532
rect 1190 528 5472 532
rect 849 520 1482 524
rect 1486 520 5472 524
rect 849 512 1994 516
rect 1998 512 5472 516
rect 849 504 2918 508
rect 2922 504 5472 508
rect 849 496 3430 500
rect 3434 496 5472 500
rect 849 488 3942 492
rect 3946 488 5472 492
rect 849 480 4454 484
rect 4458 480 5472 484
rect 849 472 4966 476
rect 4970 472 5472 476
rect 26 400 30 404
rect 849 392 1466 396
rect 1470 392 5472 396
rect 849 384 1762 388
rect 1766 384 5472 388
rect 849 376 2506 380
rect 2510 376 5472 380
rect 849 368 3018 372
rect 3022 368 5472 372
rect 849 360 3530 364
rect 3534 360 5472 364
rect 849 352 4042 356
rect 4046 352 5472 356
rect 849 344 4554 348
rect 4558 344 5472 348
rect 849 336 5066 340
rect 5070 336 5472 340
rect 26 264 30 268
rect 849 256 1746 260
rect 1750 256 5472 260
rect 849 248 2274 252
rect 2278 248 5472 252
rect 849 240 2786 244
rect 2790 240 5472 244
rect 849 232 3298 236
rect 3302 232 5472 236
rect 849 224 3810 228
rect 3814 224 5472 228
rect 849 216 4322 220
rect 4326 216 5472 220
rect 849 208 4834 212
rect 4838 208 5472 212
rect 849 200 5346 204
rect 5350 200 5472 204
rect 26 128 30 132
rect 849 120 2258 124
rect 2262 120 5472 124
rect 849 112 2770 116
rect 2774 112 5472 116
rect 849 104 3282 108
rect 3286 104 5472 108
rect 849 96 3794 100
rect 3798 96 5472 100
rect 849 88 4306 92
rect 4310 88 5472 92
rect 849 80 4818 84
rect 4822 80 5472 84
rect 849 72 5330 76
rect 5334 72 5472 76
rect 849 64 5466 68
rect 5470 64 5472 68
rect 320 56 339 60
rect 26 -8 30 -4
rect 343 -59 346 -55
rect 1864 -59 2414 -55
rect 328 -123 344 -119
rect 1863 -123 2422 -119
rect 874 -196 1870 -192
rect 1154 -211 1878 -207
rect 1434 -227 1886 -223
rect 1718 -243 1894 -239
rect 1862 -251 1982 -247
rect 2376 -283 2414 -279
rect 2418 -283 2926 -279
rect 2376 -347 2422 -343
rect 2426 -347 2934 -343
rect 598 -403 856 -399
rect 1386 -419 2382 -415
rect 1666 -434 2390 -430
rect 1950 -450 2398 -446
rect 2226 -466 2406 -462
rect 2374 -474 2494 -470
rect 2888 -506 2926 -502
rect 2930 -506 3438 -502
rect 2888 -570 2934 -566
rect 2938 -570 3446 -566
rect 1110 -626 1368 -622
rect 1898 -642 2894 -638
rect 2182 -657 2902 -653
rect 2458 -673 2910 -669
rect 2738 -689 2918 -685
rect 2886 -697 3006 -693
rect 3400 -729 3438 -725
rect 3442 -729 3950 -725
rect 3400 -793 3446 -789
rect 3450 -793 3958 -789
rect 1622 -849 1880 -845
rect 2414 -865 3406 -861
rect 2690 -880 3414 -876
rect 2970 -896 3422 -892
rect 3250 -912 3430 -908
rect 3398 -920 3518 -916
rect 3912 -952 3950 -948
rect 3954 -952 4462 -948
rect 3912 -1016 3958 -1012
rect 3962 -1016 4470 -1012
rect 2134 -1072 2392 -1068
rect 2922 -1088 3918 -1084
rect 298 -1101 332 -1097
rect 3202 -1103 3926 -1099
rect 314 -1109 340 -1105
rect 3482 -1119 3934 -1115
rect 3762 -1135 3942 -1131
rect 3910 -1143 4026 -1139
rect 4424 -1175 4462 -1171
rect 4466 -1175 4974 -1171
rect 4424 -1239 4470 -1235
rect 4474 -1239 4982 -1235
rect 2646 -1295 2904 -1291
rect 3434 -1311 4430 -1307
rect 3714 -1326 4438 -1322
rect 3994 -1342 4446 -1338
rect 4278 -1358 4454 -1354
rect 4422 -1366 4542 -1362
rect 4936 -1398 4974 -1394
rect 4978 -1398 5451 -1394
rect 4936 -1462 4982 -1458
rect 4986 -1462 5458 -1458
rect 3158 -1518 3416 -1514
rect 3946 -1534 4942 -1530
rect 4226 -1549 4950 -1545
rect 4510 -1565 4958 -1561
rect 4786 -1581 4966 -1577
rect 4934 -1589 5054 -1585
rect 3670 -1605 5074 -1601
rect 572 -1621 576 -1617
rect 856 -1621 1088 -1617
rect 1368 -1621 1600 -1617
rect 1880 -1621 2112 -1617
rect 2392 -1621 2624 -1617
rect 2904 -1621 3136 -1617
rect 3415 -1621 3649 -1617
rect 5448 -1621 5451 -1617
rect 572 -1685 576 -1681
rect 856 -1685 1088 -1681
rect 1368 -1685 1600 -1681
rect 1880 -1685 2112 -1681
rect 2392 -1685 2624 -1681
rect 2904 -1685 3136 -1681
rect 3415 -1685 3649 -1681
rect 5448 -1685 5458 -1681
rect 572 -1741 576 -1737
rect 856 -1741 1088 -1737
rect 1368 -1741 1600 -1737
rect 1880 -1741 2112 -1737
rect 2392 -1741 2624 -1737
rect 2904 -1741 3136 -1737
rect 3415 -1741 3649 -1737
<< m2contact >>
rect 332 1072 336 1076
rect 362 1064 366 1068
rect 1870 1056 1874 1060
rect 2382 1048 2386 1052
rect 2894 1040 2898 1044
rect 3406 1032 3410 1036
rect 3918 1024 3922 1028
rect 5074 1016 5078 1020
rect 2 976 6 980
rect 42 976 46 980
rect 82 976 86 980
rect 122 976 126 980
rect 162 976 166 980
rect 202 976 206 980
rect 242 976 246 980
rect 282 976 286 980
rect 346 936 350 940
rect 642 928 646 932
rect 1878 920 1882 924
rect 2390 912 2394 916
rect 2902 904 2906 908
rect 3414 896 3418 900
rect 4430 888 4434 892
rect 4942 880 4946 884
rect 626 800 630 804
rect 922 792 926 796
rect 1886 784 1890 788
rect 2398 776 2402 780
rect 2910 768 2914 772
rect 3926 760 3930 764
rect 4438 752 4442 756
rect 4950 744 4954 748
rect 906 664 910 668
rect 1202 656 1206 660
rect 1894 648 1898 652
rect 2406 640 2410 644
rect 3422 632 3426 636
rect 3934 624 3938 628
rect 4446 616 4450 620
rect 4958 608 4962 612
rect 1186 528 1190 532
rect 1482 520 1486 524
rect 1994 512 1998 516
rect 2918 504 2922 508
rect 3430 496 3434 500
rect 3942 488 3946 492
rect 4454 480 4458 484
rect 4966 472 4970 476
rect 1466 392 1470 396
rect 1762 384 1766 388
rect 2506 376 2510 380
rect 3018 368 3022 372
rect 3530 360 3534 364
rect 4042 352 4046 356
rect 4554 344 4558 348
rect 5066 336 5070 340
rect 1746 256 1750 260
rect 2274 248 2278 252
rect 2786 240 2790 244
rect 3298 232 3302 236
rect 3810 224 3814 228
rect 4322 216 4326 220
rect 4834 208 4838 212
rect 5346 200 5350 204
rect 2258 120 2262 124
rect 2770 112 2774 116
rect 3282 104 3286 108
rect 3794 96 3798 100
rect 4306 88 4310 92
rect 4818 80 4822 84
rect 5330 72 5334 76
rect 5466 64 5470 68
rect 339 56 343 60
rect 339 -59 343 -55
rect 2414 -59 2418 -55
rect 324 -123 328 -119
rect 2422 -123 2426 -119
rect 340 -179 344 -175
rect 1870 -196 1874 -192
rect 1878 -211 1882 -207
rect 1886 -227 1890 -223
rect 1714 -243 1718 -239
rect 1894 -243 1898 -239
rect 1858 -251 1862 -247
rect 2414 -283 2418 -279
rect 2926 -283 2930 -279
rect 2422 -347 2426 -343
rect 2934 -347 2938 -343
rect 594 -403 598 -399
rect 2382 -419 2386 -415
rect 2390 -434 2394 -430
rect 2398 -450 2402 -446
rect 2406 -466 2410 -462
rect 2370 -474 2374 -470
rect 2926 -506 2930 -502
rect 3438 -506 3442 -502
rect 2934 -570 2938 -566
rect 3446 -570 3450 -566
rect 1106 -626 1110 -622
rect 2894 -642 2898 -638
rect 2902 -657 2906 -653
rect 2910 -673 2914 -669
rect 2918 -689 2922 -685
rect 2882 -697 2886 -693
rect 3438 -729 3442 -725
rect 3950 -729 3954 -725
rect 3446 -793 3450 -789
rect 3958 -793 3962 -789
rect 1618 -849 1622 -845
rect 2410 -865 2414 -861
rect 3406 -865 3410 -861
rect 3414 -880 3418 -876
rect 3422 -896 3426 -892
rect 3430 -912 3434 -908
rect 3394 -920 3398 -916
rect 3950 -952 3954 -948
rect 4462 -952 4466 -948
rect 3958 -1016 3962 -1012
rect 4470 -1016 4474 -1012
rect 2130 -1072 2134 -1068
rect 3918 -1088 3922 -1084
rect 294 -1101 298 -1097
rect 332 -1101 336 -1097
rect 3926 -1103 3930 -1099
rect 310 -1109 314 -1105
rect 340 -1109 344 -1105
rect 3934 -1119 3938 -1115
rect 3942 -1135 3946 -1131
rect 3906 -1143 3910 -1139
rect 4462 -1175 4466 -1171
rect 4974 -1175 4978 -1171
rect 4470 -1239 4474 -1235
rect 4982 -1239 4986 -1235
rect 2642 -1295 2646 -1291
rect 4430 -1311 4434 -1307
rect 4438 -1326 4442 -1322
rect 4446 -1342 4450 -1338
rect 4454 -1358 4458 -1354
rect 4418 -1366 4422 -1362
rect 4974 -1398 4978 -1394
rect 5451 -1398 5455 -1394
rect 4982 -1462 4986 -1458
rect 5458 -1462 5462 -1458
rect 3154 -1518 3158 -1514
rect 4942 -1534 4946 -1530
rect 4950 -1549 4954 -1545
rect 4958 -1565 4962 -1561
rect 4966 -1581 4970 -1577
rect 4930 -1589 4934 -1585
rect 3666 -1605 3670 -1601
rect 5074 -1605 5078 -1601
rect 5451 -1621 5455 -1617
rect 526 -1661 530 -1657
rect 810 -1661 814 -1657
rect 1322 -1661 1326 -1657
rect 1834 -1661 1838 -1657
rect 2346 -1661 2350 -1657
rect 2858 -1661 2862 -1657
rect 3370 -1661 3374 -1657
rect 3882 -1661 3886 -1657
rect 4162 -1661 4166 -1657
rect 4442 -1661 4446 -1657
rect 4722 -1661 4726 -1657
rect 5002 -1661 5006 -1657
rect 5458 -1685 5462 -1681
rect 292 -1741 296 -1737
rect 5466 -1784 5470 -1780
<< metal2 >>
rect 324 -119 328 0
rect 332 -1097 336 1072
rect 339 -55 343 56
rect 346 14 350 936
rect 362 16 366 1064
rect 626 25 630 800
rect 642 16 646 928
rect 922 796 926 800
rect 906 9 910 664
rect 922 1 926 792
rect 1186 -7 1190 528
rect 1202 -15 1206 656
rect 1466 -23 1470 392
rect 1482 -31 1486 520
rect 1746 -39 1750 256
rect 1762 -47 1766 384
rect 294 -1645 298 -1101
rect 340 -1105 344 -179
rect 1870 -192 1874 1056
rect 1878 -207 1882 920
rect 310 -1645 314 -1109
rect 578 -1649 582 -234
rect 858 -267 862 -233
rect 1138 -283 1142 -226
rect 1418 -299 1422 -224
rect 1698 -315 1702 -219
rect 1858 -247 1862 -222
rect 1886 -223 1890 784
rect 1894 -239 1898 648
rect 1994 -259 1998 512
rect 2258 -263 2262 120
rect 2274 -271 2278 248
rect 594 -1645 598 -403
rect 2382 -415 2386 1048
rect 2390 -430 2394 912
rect 2210 -454 2214 -441
rect 2398 -446 2402 776
rect 1090 -1645 1094 -458
rect 2370 -470 2374 -446
rect 2406 -462 2410 640
rect 2414 -279 2418 -59
rect 2422 -343 2426 -123
rect 2506 -478 2510 376
rect 2770 -486 2774 112
rect 2786 -494 2790 240
rect 1106 -1645 1110 -626
rect 2894 -638 2898 1040
rect 2902 -653 2906 904
rect 2910 -669 2914 768
rect 2722 -681 2726 -669
rect 1602 -1645 1606 -681
rect 2882 -693 2886 -669
rect 2918 -685 2922 504
rect 2926 -502 2930 -283
rect 2934 -566 2938 -347
rect 3018 -705 3022 368
rect 3282 -709 3286 104
rect 3298 -717 3302 232
rect 1618 -1645 1622 -849
rect 3406 -861 3410 1032
rect 3414 -876 3418 896
rect 3422 -892 3426 632
rect 3234 -904 3238 -892
rect 2114 -1646 2118 -904
rect 3394 -916 3398 -892
rect 3430 -908 3434 496
rect 3438 -725 3442 -506
rect 3446 -789 3450 -570
rect 3530 -924 3534 360
rect 3794 -932 3798 96
rect 3810 -940 3814 224
rect 2130 -1645 2134 -1072
rect 3918 -1084 3922 1024
rect 3926 -1099 3930 760
rect 3934 -1115 3938 624
rect 3746 -1123 3750 -1115
rect 2626 -1645 2630 -1127
rect 3906 -1139 3910 -1115
rect 3942 -1131 3946 488
rect 3950 -948 3954 -729
rect 3958 -1012 3962 -793
rect 4042 -1147 4046 352
rect 4306 -1155 4310 88
rect 4322 -1163 4326 216
rect 2642 -1645 2646 -1295
rect 4430 -1307 4434 888
rect 4438 -1322 4442 752
rect 4446 -1338 4450 616
rect 4258 -1346 4262 -1338
rect 3138 -1665 3142 -1350
rect 4418 -1362 4422 -1338
rect 4454 -1354 4458 480
rect 4462 -1171 4466 -952
rect 4470 -1235 4474 -1016
rect 4554 -1370 4558 344
rect 4818 -1378 4822 80
rect 4834 -1386 4838 208
rect 3154 -1665 3158 -1518
rect 4942 -1530 4946 880
rect 4950 -1545 4954 744
rect 4958 -1561 4962 608
rect 4770 -1573 4774 -1561
rect 3650 -1645 3654 -1573
rect 4930 -1585 4934 -1561
rect 4966 -1577 4970 472
rect 4974 -1394 4978 -1175
rect 4982 -1458 4986 -1239
rect 5066 -1597 5070 336
rect 5074 -1601 5078 1016
rect 5330 -1605 5334 72
rect 3666 -1649 3670 -1605
rect 5346 -1609 5350 200
rect 5451 -1617 5455 -1398
rect 5458 -1681 5462 -1462
rect 5466 -1780 5470 64
rect 4162 -1828 4166 -1796
rect 4442 -1820 4446 -1796
rect 4722 -1812 4726 -1792
rect 5002 -1804 5006 -1788
rect 5282 -1796 5286 -1784
rect 5442 -1788 5446 -1784
use Add5  Add5_0
timestamp 1714258260
transform 1 0 624 0 1 -123
box -284 -111 1242 163
use Add5  Add5_1
timestamp 1714258260
transform 1 0 1136 0 1 -347
box -284 -111 1242 163
use Add5  Add5_2
timestamp 1714258260
transform 1 0 1648 0 1 -570
box -284 -111 1242 163
use Add5  Add5_3
timestamp 1714258260
transform 1 0 2160 0 1 -793
box -284 -111 1242 163
use Add5  Add5_4
timestamp 1714258260
transform 1 0 2672 0 1 -1016
box -284 -111 1242 163
use Add5  Add5_5
timestamp 1714258260
transform 1 0 3184 0 1 -1239
box -284 -111 1242 163
use Add5  Add5_6
timestamp 1714258260
transform 1 0 3696 0 1 -1462
box -284 -111 1242 163
use Add5  Add5_7
timestamp 1714258260
transform 1 0 4208 0 1 -1685
box -284 -111 1242 163
use M_FA  M_FA_0
timestamp 1714172470
transform 1 0 3648 0 1 -1685
box -4 -56 284 71
use M_FA  M_FA_1
timestamp 1714172470
transform 1 0 3136 0 1 -1685
box -4 -56 284 71
use M_FA  M_FA_2
timestamp 1714172470
transform 1 0 2624 0 1 -1685
box -4 -56 284 71
use M_FA  M_FA_3
timestamp 1714172470
transform 1 0 2112 0 1 -1685
box -4 -56 284 71
use M_FA  M_FA_4
timestamp 1714172470
transform 1 0 1600 0 1 -1685
box -4 -56 284 71
use M_FA  M_FA_5
timestamp 1714172470
transform 1 0 1088 0 1 -1685
box -4 -56 284 71
use M_FA  M_FA_6
timestamp 1714172470
transform 1 0 576 0 1 -1685
box -4 -56 284 71
use M_FA  M_FA_7
timestamp 1714172470
transform 1 0 292 0 1 -1685
box -4 -56 284 71
use Partial  Partial_0
timestamp 1714342102
transform 1 0 0 0 1 952
box -8 -960 892 124
<< labels >>
rlabel m2contact 5468 -1782 5468 -1782 7 q0
rlabel metal1 1 954 1 954 1 VSS
rlabel m2contact 4 978 4 978 1 A7
rlabel m2contact 44 978 44 978 1 A6
rlabel m2contact 84 978 84 978 1 A5
rlabel m2contact 124 978 124 978 1 A4
rlabel m2contact 164 978 164 978 1 A3
rlabel m2contact 204 978 204 978 1 A2
rlabel m2contact 244 978 244 978 1 A1
rlabel m2contact 284 978 284 978 1 A0
rlabel metal1 28 -6 28 -6 1 M0
rlabel metal1 28 130 28 130 1 M1
rlabel metal1 28 266 28 266 1 M2
rlabel metal1 28 402 28 402 1 M3
rlabel metal1 28 538 28 538 1 M4
rlabel metal1 28 674 28 674 1 M5
rlabel metal1 28 810 28 810 1 M6
rlabel metal1 28 946 28 946 1 M7
rlabel metal2 1698 -235 1702 -231 1 q4_A
rlabel metal2 5444 -1786 5444 -1786 1 q1
rlabel metal2 5284 -1786 5284 -1786 1 q2
rlabel m2contact 5004 -1659 5004 -1659 1 q3
rlabel m2contact 4724 -1659 4724 -1659 1 q4
rlabel m2contact 4444 -1659 4444 -1659 1 q5
rlabel m2contact 4164 -1659 4164 -1659 1 q6
rlabel m2contact 3884 -1659 3884 -1659 1 q7
rlabel m2contact 3372 -1659 3372 -1659 1 q8
rlabel m2contact 2860 -1659 2860 -1659 1 q9
rlabel m2contact 2348 -1659 2348 -1659 1 q10
rlabel m2contact 1836 -1659 1836 -1659 1 q11
rlabel m2contact 1324 -1659 1324 -1659 1 q12
rlabel m2contact 812 -1659 812 -1659 1 q13
rlabel m2contact 528 -1659 528 -1659 1 q14
rlabel m2contact 294 -1739 294 -1739 1 q15
rlabel metal1 -2 1010 -2 1010 1 VDD
<< end >>
