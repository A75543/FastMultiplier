magic
tech scmos
timestamp 1715208163
<< nwell >>
rect 165 3792 171 3794
rect 2834 1159 2843 1163
rect 1869 275 1871 279
<< polycontact >>
rect 1340 4278 1344 4282
rect 1356 4278 1360 4282
rect 1372 4278 1376 4282
rect 1388 4278 1392 4282
rect 1404 4278 1408 4282
rect 1420 4278 1424 4282
rect 1436 4278 1440 4282
rect 1452 4278 1456 4282
<< metal1 >>
rect 158 4034 164 4038
rect 174 4034 180 4038
rect 190 4034 197 4038
rect 246 3978 250 3982
rect 314 3978 365 3982
rect 426 3978 477 3982
rect 538 3978 589 3982
rect 650 3978 701 3982
rect 762 3978 813 3982
rect 874 3978 925 3982
rect 986 3978 1037 3982
rect 1098 3978 1149 3982
rect 168 3914 172 3918
rect 260 3914 278 3918
rect 284 3914 294 3918
rect 247 3849 251 3853
rect 166 3788 170 3792
rect 260 3788 270 3792
rect 276 3788 286 3792
rect 300 3788 308 3792
rect 1247 3788 1251 3792
rect 108 3724 116 3745
rect 207 3731 212 3736
rect 3626 1828 3632 1832
rect 3642 1828 3658 1832
rect 3664 1828 3669 1832
rect 3730 1828 3736 1832
rect 3746 1828 3752 1832
rect 3762 1828 3776 1832
rect 3842 1828 3856 1832
rect 3866 1828 3880 1832
rect 2162 1159 2213 1163
rect 2274 1159 2312 1163
rect 2386 1159 2395 1163
rect 2399 1159 2435 1163
rect 2498 1159 2515 1163
rect 2519 1159 2549 1163
rect 2610 1159 2661 1163
rect 2722 1159 2773 1163
rect 2871 1159 2883 1163
rect 2951 1159 2963 1163
rect 2967 1159 2987 1163
rect 2991 1159 2997 1163
rect 3058 1159 3067 1163
rect 3071 1159 3091 1163
rect 3095 1159 3109 1163
rect 3170 1159 3221 1163
rect 3282 1159 3333 1163
rect 3399 1159 3419 1163
rect 3423 1159 3445 1163
rect 3506 1159 3515 1163
rect 3519 1159 3539 1163
rect 3618 1159 3669 1163
rect 3730 1159 3781 1163
rect 3842 1159 3848 1163
rect 3858 1159 3864 1163
rect 3874 1159 3891 1163
rect 3975 1159 3987 1163
rect 3991 1159 4005 1163
rect 4066 1159 4091 1163
rect 4095 1159 4115 1163
rect 4290 1159 4341 1163
rect 4407 1159 4419 1163
rect 4423 1159 4443 1163
rect 4447 1159 4453 1163
rect 4514 1159 4523 1163
rect 4527 1159 4539 1163
rect 4543 1159 4563 1163
rect 4631 1159 4677 1163
rect 4738 1159 4789 1163
rect 4850 1159 4872 1163
rect 4882 1159 4888 1163
rect 4962 1159 4995 1163
rect 4999 1159 5011 1163
rect 5079 1159 5115 1163
rect 5119 1159 5125 1163
rect 5186 1159 5195 1163
rect 5199 1159 5211 1163
rect 5215 1159 5235 1163
rect 5298 1159 5315 1163
rect 5319 1159 5331 1163
rect 5335 1159 5349 1163
rect 5410 1159 5419 1163
rect 5423 1159 5432 1163
rect 5442 1159 5448 1163
rect 5522 1159 5555 1163
rect 5559 1159 5571 1163
rect 5639 1159 5675 1163
rect 5679 1159 5683 1163
rect 5746 1159 5755 1163
rect 5760 1159 5771 1163
rect 5775 1159 5795 1163
rect 5858 1159 5875 1163
rect 5879 1159 5891 1163
rect 5896 1159 5909 1163
rect 5970 1159 5979 1163
rect 5984 1159 5992 1163
rect 6002 1159 6008 1163
rect 6082 1159 6115 1163
rect 6199 1159 6235 1163
rect 6306 1159 6315 1163
rect 6320 1159 6331 1163
rect 6335 1159 6355 1163
rect 6418 1159 6435 1163
rect 6439 1159 6451 1163
rect 6455 1159 6469 1163
rect 6530 1159 6539 1163
rect 1826 275 1833 279
rect 1837 275 1869 279
rect 1938 275 1953 279
rect 1957 275 1989 279
rect 2053 275 2073 279
rect 2077 275 2101 279
rect 2162 275 2168 279
rect 2172 275 2192 279
rect 2196 275 2213 279
rect 2276 275 2288 279
rect 2292 275 2312 279
rect 2316 275 2325 279
rect 2386 275 2392 279
rect 2396 275 2408 279
rect 2412 275 2432 279
rect 2498 275 2512 279
rect 2516 275 2528 279
rect 2532 275 2549 279
rect 2612 275 2632 279
rect 2636 275 2648 279
rect 2652 275 2661 279
rect 1882 211 1886 215
rect 1997 211 1999 215
rect 2001 211 2006 215
rect 2239 211 2245 215
rect 2359 211 2365 215
rect 2479 211 2485 215
rect 2599 211 2605 215
rect 2711 211 2717 215
rect 2778 211 2829 215
rect 2728 149 2734 153
rect 1817 93 1821 97
rect 2112 93 2118 97
rect 2196 93 2200 97
rect 2386 93 2390 97
rect 2670 93 2674 97
rect 2685 93 2689 97
rect 2790 93 2800 97
rect 1788 89 1792 93
rect 1925 89 1929 93
rect 2005 89 2009 93
<< m2contact >>
rect 1227 4032 1231 4036
rect 119 3998 123 4002
rect 135 3998 139 4002
rect 151 3998 155 4002
rect 167 3998 171 4002
rect 183 3998 187 4002
rect 199 3998 203 4002
rect 215 3998 219 4002
rect 231 3998 235 4002
rect 116 3982 120 3986
rect 145 3788 149 3792
rect 16 3732 20 3736
rect 340 3731 350 3736
rect 1881 557 1885 561
rect 2017 557 2021 561
rect 2153 557 2157 561
rect 2289 557 2293 561
rect 2425 557 2429 561
rect 2561 557 2565 561
rect 2697 557 2701 561
rect 2833 557 2837 561
rect 1881 105 1885 109
rect 2017 105 2021 109
rect 2153 105 2157 109
rect 2289 105 2293 109
rect 2425 105 2429 109
rect 2561 105 2565 109
rect 2697 105 2701 109
rect 2833 105 2837 109
<< metal2 >>
rect 145 3792 146 3793
rect 149 3788 150 3792
<< m3contact >>
rect 158 4034 164 4038
rect 174 4034 180 4038
rect 190 4034 197 4038
rect 116 3986 121 3991
rect 246 3978 251 3984
rect 314 3978 365 3982
rect 426 3978 477 3982
rect 538 3978 589 3982
rect 650 3978 701 3982
rect 762 3978 813 3982
rect 874 3978 925 3982
rect 986 3978 1037 3982
rect 1098 3978 1149 3982
rect 167 3913 173 3919
rect 260 3914 278 3918
rect 284 3914 294 3918
rect 247 3848 252 3853
rect 146 3792 151 3797
rect 165 3788 171 3792
rect 260 3788 270 3792
rect 276 3788 286 3792
rect 300 3788 308 3792
rect 1247 3788 1251 3792
rect 15 3727 20 3732
rect 108 3724 116 3745
rect 207 3730 213 3736
rect 3626 1828 3632 1832
rect 3642 1828 3658 1832
rect 3664 1828 3669 1832
rect 3730 1828 3736 1832
rect 3746 1828 3752 1832
rect 3762 1828 3776 1832
rect 3842 1828 3856 1832
rect 3866 1828 3880 1832
rect 2162 1159 2213 1163
rect 2274 1159 2312 1163
rect 2386 1159 2395 1163
rect 2399 1159 2435 1163
rect 2498 1159 2515 1163
rect 2519 1159 2549 1163
rect 2610 1159 2661 1163
rect 2722 1159 2773 1163
rect 2871 1159 2883 1163
rect 2951 1159 2963 1163
rect 2967 1159 2987 1163
rect 2991 1159 2997 1163
rect 3058 1159 3067 1163
rect 3071 1159 3091 1163
rect 3095 1159 3109 1163
rect 3170 1159 3221 1163
rect 3282 1159 3333 1163
rect 3399 1159 3419 1163
rect 3423 1159 3445 1163
rect 3506 1159 3515 1163
rect 3519 1159 3539 1163
rect 3618 1159 3669 1163
rect 3730 1159 3781 1163
rect 3842 1159 3848 1163
rect 3858 1159 3864 1163
rect 3874 1159 3891 1163
rect 3956 1159 3971 1163
rect 3975 1159 3987 1163
rect 3991 1159 4005 1163
rect 4066 1159 4091 1163
rect 4095 1159 4115 1163
rect 4178 1159 4229 1163
rect 4290 1159 4341 1163
rect 4407 1159 4419 1163
rect 4423 1159 4443 1163
rect 4447 1159 4453 1163
rect 4514 1159 4523 1163
rect 4527 1159 4539 1163
rect 4543 1159 4563 1163
rect 4631 1159 4677 1163
rect 4738 1159 4789 1163
rect 4850 1159 4872 1163
rect 4882 1159 4888 1163
rect 4962 1159 4995 1163
rect 4999 1159 5011 1163
rect 5079 1159 5115 1163
rect 5119 1159 5125 1163
rect 5186 1159 5195 1163
rect 5199 1159 5211 1163
rect 5215 1159 5235 1163
rect 5298 1159 5315 1163
rect 5319 1159 5331 1163
rect 5335 1159 5349 1163
rect 5410 1159 5419 1163
rect 5423 1159 5432 1163
rect 5442 1159 5448 1163
rect 5522 1159 5555 1163
rect 5559 1159 5571 1163
rect 5639 1159 5675 1163
rect 5679 1159 5683 1163
rect 5746 1159 5755 1163
rect 5760 1159 5771 1163
rect 5775 1159 5795 1163
rect 5858 1159 5875 1163
rect 5879 1159 5891 1163
rect 5896 1159 5909 1163
rect 5970 1159 5979 1163
rect 5984 1159 5992 1163
rect 6002 1159 6008 1163
rect 6082 1159 6115 1163
rect 6119 1159 6131 1163
rect 6199 1159 6235 1163
rect 6306 1159 6315 1163
rect 6320 1159 6331 1163
rect 6335 1159 6355 1163
rect 6418 1159 6435 1163
rect 6439 1159 6451 1163
rect 6455 1159 6469 1163
rect 6530 1159 6539 1163
rect 6642 1159 6673 1163
rect 1743 605 1748 610
rect 1826 275 1833 279
rect 1837 275 1869 279
rect 1938 275 1953 279
rect 1957 275 1989 279
rect 2053 275 2073 279
rect 2077 275 2101 279
rect 2162 275 2168 279
rect 2172 275 2192 279
rect 2196 275 2213 279
rect 2276 275 2288 279
rect 2292 275 2312 279
rect 2316 275 2325 279
rect 2386 275 2392 279
rect 2396 275 2408 279
rect 2412 275 2432 279
rect 2498 275 2512 279
rect 2516 275 2528 279
rect 2532 275 2549 279
rect 2612 275 2632 279
rect 2636 275 2648 279
rect 2652 275 2661 279
rect 1882 211 1886 215
rect 2001 211 2006 215
rect 2239 211 2245 215
rect 2359 211 2365 215
rect 2479 211 2485 215
rect 2599 211 2605 215
rect 2711 211 2717 215
rect 2778 211 2829 215
rect 2728 149 2734 153
rect 2112 93 2118 97
rect 2196 93 2200 97
rect 2386 93 2390 97
rect 2670 93 2674 97
rect 2685 93 2689 97
rect 2790 93 2800 97
rect 1788 89 1792 93
rect 1925 89 1929 93
rect 2005 89 2009 93
<< metal3 >>
rect -23 4320 6750 4332
rect -23 3732 30 4320
rect -23 3727 15 3732
rect 20 3727 30 3732
rect -23 9 30 3727
rect 33 6 86 4317
rect 89 3991 142 4320
rect 89 3986 116 3991
rect 121 3986 142 3991
rect 89 3745 142 3986
rect 89 3724 108 3745
rect 116 3724 142 3745
rect 89 9 142 3724
rect 145 4038 198 4317
rect 145 4034 158 4038
rect 164 4034 174 4038
rect 180 4034 190 4038
rect 197 4034 198 4038
rect 145 3919 198 4034
rect 145 3913 167 3919
rect 173 3913 198 3919
rect 145 3797 198 3913
rect 145 3792 146 3797
rect 151 3792 198 3797
rect 145 3788 165 3792
rect 171 3788 198 3792
rect 145 6 198 3788
rect 201 3984 254 4320
rect 201 3978 246 3984
rect 251 3978 254 3984
rect 201 3853 254 3978
rect 201 3848 247 3853
rect 252 3848 254 3853
rect 201 3736 254 3848
rect 201 3730 207 3736
rect 213 3730 254 3736
rect 201 9 254 3730
rect 257 3918 310 4317
rect 257 3914 260 3918
rect 278 3914 284 3918
rect 294 3914 310 3918
rect 257 3792 310 3914
rect 257 3788 260 3792
rect 270 3788 276 3792
rect 286 3788 300 3792
rect 308 3788 310 3792
rect 257 6 310 3788
rect 313 3982 366 4320
rect 313 3978 314 3982
rect 365 3978 366 3982
rect 313 9 366 3978
rect 369 6 422 4317
rect 425 3982 478 4320
rect 425 3978 426 3982
rect 477 3978 478 3982
rect 425 9 478 3978
rect 481 6 534 4317
rect 537 3982 590 4320
rect 537 3978 538 3982
rect 589 3978 590 3982
rect 537 9 590 3978
rect 593 6 646 4317
rect 649 3982 702 4320
rect 649 3978 650 3982
rect 701 3978 702 3982
rect 649 9 702 3978
rect 705 6 758 4317
rect 761 3982 814 4320
rect 761 3978 762 3982
rect 813 3978 814 3982
rect 761 9 814 3978
rect 817 6 870 4317
rect 873 3982 926 4320
rect 873 3978 874 3982
rect 925 3978 926 3982
rect 873 9 926 3978
rect 929 6 982 4317
rect 985 3982 1038 4320
rect 985 3978 986 3982
rect 1037 3978 1038 3982
rect 985 9 1038 3978
rect 1041 6 1094 4317
rect 1097 3982 1150 4320
rect 1097 3978 1098 3982
rect 1149 3978 1150 3982
rect 1097 9 1150 3978
rect 1153 6 1206 4317
rect 1209 3792 1262 4320
rect 1209 3788 1247 3792
rect 1251 3788 1262 3792
rect 1209 9 1262 3788
rect 1265 6 1318 4317
rect 1321 9 1374 4320
rect 1377 4282 1430 4317
rect 1377 4278 1388 4282
rect 1392 4278 1430 4282
rect 1377 6 1430 4278
rect 1433 9 1486 4320
rect 1489 6 1542 4317
rect 1545 9 1598 4320
rect 1601 6 1654 4317
rect 1657 9 1710 4320
rect 1713 610 1766 4317
rect 1713 605 1743 610
rect 1748 605 1766 610
rect 1713 6 1766 605
rect 1769 93 1822 4320
rect 1769 89 1788 93
rect 1792 89 1822 93
rect 1769 9 1822 89
rect 1825 279 1878 4317
rect 1825 275 1826 279
rect 1833 275 1837 279
rect 1869 275 1878 279
rect 1825 6 1878 275
rect 1881 215 1934 4320
rect 1881 211 1882 215
rect 1886 211 1934 215
rect 1881 93 1934 211
rect 1881 89 1925 93
rect 1929 89 1934 93
rect 1881 9 1934 89
rect 1937 279 1990 4317
rect 1937 275 1938 279
rect 1953 275 1957 279
rect 1989 275 1990 279
rect 1937 6 1990 275
rect 1993 215 2046 4320
rect 1993 211 2001 215
rect 2006 211 2046 215
rect 1993 93 2046 211
rect 1993 89 2005 93
rect 2009 89 2046 93
rect 1993 9 2046 89
rect 2049 279 2102 4316
rect 2049 275 2053 279
rect 2073 275 2077 279
rect 2101 275 2102 279
rect 2049 6 2102 275
rect 2105 97 2158 4320
rect 2105 93 2112 97
rect 2118 93 2158 97
rect 2105 9 2158 93
rect 2161 1163 2214 4317
rect 2161 1159 2162 1163
rect 2213 1159 2214 1163
rect 2161 279 2214 1159
rect 2161 275 2162 279
rect 2168 275 2172 279
rect 2192 275 2196 279
rect 2213 275 2214 279
rect 2161 97 2214 275
rect 2161 93 2196 97
rect 2200 93 2214 97
rect 2161 6 2214 93
rect 2217 215 2270 4320
rect 2217 211 2239 215
rect 2245 211 2270 215
rect 2217 9 2270 211
rect 2273 1163 2326 4317
rect 2273 1159 2274 1163
rect 2312 1159 2326 1163
rect 2273 279 2326 1159
rect 2273 275 2276 279
rect 2288 275 2292 279
rect 2312 275 2316 279
rect 2325 275 2326 279
rect 2273 6 2326 275
rect 2329 215 2382 4320
rect 2329 211 2359 215
rect 2365 211 2382 215
rect 2329 9 2382 211
rect 2385 1163 2438 4317
rect 2385 1159 2386 1163
rect 2395 1159 2399 1163
rect 2435 1159 2438 1163
rect 2385 279 2438 1159
rect 2385 275 2386 279
rect 2392 275 2396 279
rect 2408 275 2412 279
rect 2432 275 2438 279
rect 2385 97 2438 275
rect 2385 93 2386 97
rect 2390 93 2438 97
rect 2385 6 2438 93
rect 2441 215 2494 4320
rect 2441 211 2479 215
rect 2485 211 2494 215
rect 2441 9 2494 211
rect 2497 1163 2550 4317
rect 2497 1159 2498 1163
rect 2515 1159 2519 1163
rect 2549 1159 2550 1163
rect 2497 279 2550 1159
rect 2497 275 2498 279
rect 2512 275 2516 279
rect 2528 275 2532 279
rect 2549 275 2550 279
rect 2497 6 2550 275
rect 2553 215 2606 4320
rect 2553 211 2599 215
rect 2605 211 2606 215
rect 2553 9 2606 211
rect 2609 1163 2662 4317
rect 2609 1159 2610 1163
rect 2661 1159 2662 1163
rect 2609 279 2662 1159
rect 2609 275 2612 279
rect 2632 275 2636 279
rect 2648 275 2652 279
rect 2661 275 2662 279
rect 2609 6 2662 275
rect 2665 215 2718 4320
rect 2665 211 2711 215
rect 2717 211 2718 215
rect 2665 97 2718 211
rect 2665 93 2670 97
rect 2674 93 2685 97
rect 2689 93 2718 97
rect 2665 9 2718 93
rect 2721 1163 2774 4317
rect 2721 1159 2722 1163
rect 2773 1159 2774 1163
rect 2721 153 2774 1159
rect 2721 149 2728 153
rect 2734 149 2774 153
rect 2721 6 2774 149
rect 2777 215 2830 4320
rect 2777 211 2778 215
rect 2829 211 2830 215
rect 2777 97 2830 211
rect 2833 1163 2886 4317
rect 2833 1159 2871 1163
rect 2883 1159 2886 1163
rect 2833 109 2886 1159
rect 2837 105 2886 109
rect 2777 93 2790 97
rect 2800 93 2830 97
rect 2777 9 2830 93
rect 2833 6 2886 105
rect 2889 9 2942 4320
rect 2945 1163 2998 4317
rect 2945 1159 2951 1163
rect 2963 1159 2967 1163
rect 2987 1159 2991 1163
rect 2997 1159 2998 1163
rect 2945 6 2998 1159
rect 3001 9 3054 4320
rect 3057 1163 3110 4317
rect 3057 1159 3058 1163
rect 3067 1159 3071 1163
rect 3091 1159 3095 1163
rect 3109 1159 3110 1163
rect 3057 6 3110 1159
rect 3113 9 3166 4320
rect 3169 1163 3222 4317
rect 3169 1159 3170 1163
rect 3221 1159 3222 1163
rect 3169 6 3222 1159
rect 3225 9 3278 4320
rect 3281 1163 3334 4317
rect 3281 1159 3282 1163
rect 3333 1159 3334 1163
rect 3281 6 3334 1159
rect 3337 9 3390 4320
rect 3393 1163 3446 4317
rect 3393 1159 3399 1163
rect 3419 1159 3423 1163
rect 3445 1159 3446 1163
rect 3393 6 3446 1159
rect 3449 9 3502 4320
rect 3505 1163 3558 4317
rect 3505 1159 3506 1163
rect 3515 1159 3519 1163
rect 3539 1159 3558 1163
rect 3505 6 3558 1159
rect 3561 9 3614 4320
rect 3617 1832 3670 4317
rect 3617 1828 3626 1832
rect 3632 1828 3642 1832
rect 3658 1828 3664 1832
rect 3669 1828 3670 1832
rect 3617 1163 3670 1828
rect 3617 1159 3618 1163
rect 3669 1159 3670 1163
rect 3617 6 3670 1159
rect 3673 9 3726 4320
rect 3729 1832 3782 4317
rect 3729 1828 3730 1832
rect 3736 1828 3746 1832
rect 3752 1828 3762 1832
rect 3776 1828 3782 1832
rect 3729 1163 3782 1828
rect 3729 1159 3730 1163
rect 3781 1159 3782 1163
rect 3729 6 3782 1159
rect 3785 9 3838 4320
rect 3841 1832 3894 4317
rect 3841 1828 3842 1832
rect 3856 1828 3866 1832
rect 3880 1828 3894 1832
rect 3841 1163 3894 1828
rect 3841 1159 3842 1163
rect 3848 1159 3858 1163
rect 3864 1159 3874 1163
rect 3891 1159 3894 1163
rect 3841 6 3894 1159
rect 3897 9 3950 4320
rect 3953 1163 4006 4317
rect 3953 1159 3956 1163
rect 3971 1159 3975 1163
rect 3987 1159 3991 1163
rect 4005 1159 4006 1163
rect 3953 6 4006 1159
rect 4009 9 4062 4320
rect 4065 1163 4118 4317
rect 4065 1159 4066 1163
rect 4091 1159 4095 1163
rect 4115 1159 4118 1163
rect 4065 6 4118 1159
rect 4121 9 4174 4320
rect 4177 1163 4230 4317
rect 4177 1159 4178 1163
rect 4229 1159 4230 1163
rect 4177 6 4230 1159
rect 4233 9 4286 4320
rect 4289 1163 4342 4317
rect 4289 1159 4290 1163
rect 4341 1159 4342 1163
rect 4289 6 4342 1159
rect 4345 9 4398 4320
rect 4401 1163 4454 4317
rect 4401 1159 4407 1163
rect 4419 1159 4423 1163
rect 4443 1159 4447 1163
rect 4453 1159 4454 1163
rect 4401 6 4454 1159
rect 4457 9 4510 4320
rect 4513 1163 4566 4317
rect 4513 1159 4514 1163
rect 4523 1159 4527 1163
rect 4539 1159 4543 1163
rect 4563 1159 4566 1163
rect 4513 6 4566 1159
rect 4569 9 4622 4320
rect 4625 1163 4678 4317
rect 4625 1159 4631 1163
rect 4677 1159 4678 1163
rect 4625 6 4678 1159
rect 4681 9 4734 4320
rect 4737 1163 4790 4317
rect 4737 1159 4738 1163
rect 4789 1159 4790 1163
rect 4737 6 4790 1159
rect 4793 9 4846 4320
rect 4849 1163 4902 4317
rect 4849 1159 4850 1163
rect 4872 1159 4882 1163
rect 4888 1159 4902 1163
rect 4849 6 4902 1159
rect 4905 9 4958 4320
rect 4961 1163 5014 4317
rect 4961 1159 4962 1163
rect 4995 1159 4999 1163
rect 5011 1159 5014 1163
rect 4961 6 5014 1159
rect 5017 9 5070 4320
rect 5073 1163 5126 4317
rect 5073 1159 5079 1163
rect 5115 1159 5119 1163
rect 5125 1159 5126 1163
rect 5073 6 5126 1159
rect 5129 9 5182 4320
rect 5185 1163 5238 4317
rect 5185 1159 5186 1163
rect 5195 1159 5199 1163
rect 5211 1159 5215 1163
rect 5235 1159 5238 1163
rect 5185 6 5238 1159
rect 5241 9 5294 4320
rect 5297 1163 5350 4317
rect 5297 1159 5298 1163
rect 5315 1159 5319 1163
rect 5331 1159 5335 1163
rect 5349 1159 5350 1163
rect 5297 6 5350 1159
rect 5353 9 5406 4320
rect 5409 1163 5462 4317
rect 5409 1159 5410 1163
rect 5419 1159 5423 1163
rect 5432 1159 5442 1163
rect 5448 1159 5462 1163
rect 5409 6 5462 1159
rect 5465 9 5518 4320
rect 5521 1163 5574 4317
rect 5521 1159 5522 1163
rect 5555 1159 5559 1163
rect 5571 1159 5574 1163
rect 5521 6 5574 1159
rect 5577 9 5630 4320
rect 5633 1163 5686 4317
rect 5633 1159 5639 1163
rect 5675 1159 5679 1163
rect 5683 1159 5686 1163
rect 5633 6 5686 1159
rect 5689 9 5742 4320
rect 5745 1163 5798 4317
rect 5745 1159 5746 1163
rect 5755 1159 5760 1163
rect 5771 1159 5775 1163
rect 5795 1159 5798 1163
rect 5745 6 5798 1159
rect 5801 9 5854 4320
rect 5857 1163 5910 4317
rect 5857 1159 5858 1163
rect 5875 1159 5879 1163
rect 5891 1159 5896 1163
rect 5909 1159 5910 1163
rect 5857 6 5910 1159
rect 5913 9 5966 4320
rect 5969 1163 6022 4317
rect 5969 1159 5970 1163
rect 5979 1159 5984 1163
rect 5992 1159 6002 1163
rect 6008 1159 6022 1163
rect 5969 6 6022 1159
rect 6025 9 6078 4320
rect 6081 1163 6134 4317
rect 6081 1159 6082 1163
rect 6115 1159 6119 1163
rect 6131 1159 6134 1163
rect 6081 6 6134 1159
rect 6137 9 6190 4320
rect 6193 1163 6246 4317
rect 6193 1159 6199 1163
rect 6235 1159 6246 1163
rect 6193 6 6246 1159
rect 6249 9 6302 4320
rect 6305 1163 6358 4317
rect 6305 1159 6306 1163
rect 6315 1159 6320 1163
rect 6331 1159 6335 1163
rect 6355 1159 6358 1163
rect 6305 6 6358 1159
rect 6361 9 6414 4320
rect 6417 1163 6470 4317
rect 6417 1159 6418 1163
rect 6435 1159 6439 1163
rect 6451 1159 6455 1163
rect 6469 1159 6470 1163
rect 6417 6 6470 1159
rect 6473 9 6526 4320
rect 6529 1163 6582 4317
rect 6529 1159 6530 1163
rect 6539 1159 6582 1163
rect 6529 6 6582 1159
rect 6585 9 6638 4320
rect 6641 1163 6694 4317
rect 6641 1159 6642 1163
rect 6673 1159 6694 1163
rect 6641 6 6694 1159
rect 6697 9 6750 4320
rect -23 -6 6750 6
use Multiplier  Multiplier_1
timestamp 1715207069
transform 1 0 1225 0 1 4008
box -1225 -4008 5472 318
<< labels >>
rlabel m2contact 1229 4034 1229 4034 1 Sign
rlabel metal3 -23 3732 30 4326 1 VSS
rlabel metal3 -23 0 6750 6 1 VDD
rlabel m2contact 1883 559 1883 559 1 Q0
rlabel m2contact 2019 559 2019 559 1 Q1
rlabel m2contact 2155 559 2155 559 1 Q2
rlabel m2contact 2291 559 2291 559 1 Q3
rlabel m2contact 2427 559 2427 559 1 Q4
rlabel m2contact 2563 559 2563 559 1 Q5
rlabel m2contact 2699 559 2699 559 1 Q6
rlabel m2contact 2835 559 2835 559 1 Q7
rlabel m2contact 1883 107 1883 107 1 Q8
rlabel m2contact 2019 107 2019 107 1 Q9
rlabel m2contact 2155 107 2155 107 1 Q10
rlabel m2contact 2291 107 2291 107 1 Q11
rlabel m2contact 2427 107 2427 107 1 Q12
rlabel m2contact 2563 107 2563 107 1 Q13
rlabel m2contact 2699 107 2699 107 1 Q14
rlabel m2contact 2835 107 2835 107 1 Q15
rlabel polycontact 1342 4280 1342 4280 1 A0
rlabel polycontact 1358 4280 1358 4280 1 A1
rlabel polycontact 1374 4280 1374 4280 1 A2
rlabel polycontact 1390 4280 1390 4280 1 A3
rlabel polycontact 1406 4280 1406 4280 1 A4
rlabel polycontact 1422 4280 1422 4280 1 A5
rlabel polycontact 1438 4280 1438 4280 1 A6
rlabel polycontact 1454 4280 1454 4280 1 A7
rlabel m2contact 121 4000 121 4000 1 B0
rlabel m2contact 137 4000 137 4000 1 B1
rlabel m2contact 153 4000 153 4000 1 B2
rlabel m2contact 169 4000 169 4000 1 B3
rlabel m2contact 185 4000 185 4000 1 B4
rlabel m2contact 201 4000 201 4000 1 B5
rlabel m2contact 217 4000 217 4000 1 B6
rlabel m2contact 233 4000 233 4000 1 B7
<< end >>
