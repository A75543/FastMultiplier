magic
tech scmos
timestamp 1711559697
<< nwell >>
rect -4 30 44 66
<< ntransistor >>
rect 7 8 9 12
rect 15 8 17 12
rect 31 8 33 12
<< ptransistor >>
rect 7 36 9 52
rect 15 36 17 52
rect 31 36 33 52
<< ndiffusion >>
rect 6 8 7 12
rect 9 8 10 12
rect 14 8 15 12
rect 17 8 18 12
rect 30 8 31 12
rect 33 8 34 12
<< pdiffusion >>
rect 6 36 7 52
rect 9 36 15 52
rect 17 36 18 52
rect 30 36 31 52
rect 33 36 34 52
<< ndcontact >>
rect 2 8 6 12
rect 10 8 14 12
rect 18 8 22 12
rect 26 8 30 12
rect 34 8 38 12
<< pdcontact >>
rect 2 36 6 52
rect 18 36 22 52
rect 26 36 30 52
rect 34 36 38 52
<< psubstratepcontact >>
rect 2 0 6 4
rect 18 0 22 4
rect 26 0 30 4
<< nsubstratencontact >>
rect 2 56 6 60
rect 26 56 30 60
<< polysilicon >>
rect 7 52 9 54
rect 15 52 17 54
rect 31 52 33 54
rect 7 32 9 36
rect 6 28 9 32
rect 7 12 9 28
rect 15 20 17 36
rect 31 28 33 36
rect 30 24 33 28
rect 15 16 18 20
rect 15 12 17 16
rect 31 12 33 24
rect 7 6 9 8
rect 15 6 17 8
rect 31 6 33 8
<< polycontact >>
rect 2 28 6 32
rect 26 24 30 28
rect 18 16 22 20
<< metal1 >>
rect 0 56 2 60
rect 6 56 26 60
rect 30 56 40 60
rect 2 52 6 56
rect 26 52 30 56
rect 18 28 22 36
rect 10 24 26 28
rect 10 12 14 24
rect 34 12 38 36
rect 2 4 6 8
rect 18 4 22 8
rect 26 4 30 8
rect 0 0 2 4
rect 6 0 18 4
rect 22 0 26 4
rect 30 0 40 4
<< labels >>
rlabel polycontact 20 18 20 18 7 B
rlabel psubstratepcontact 4 2 4 2 2 VSS
rlabel psubstratepcontact 20 2 20 2 8 VSS
rlabel psubstratepcontact 28 2 28 2 1 VSS
rlabel nsubstratencontact 4 58 4 58 4 VDD
rlabel polycontact 4 30 4 30 3 A
rlabel metal1 36 26 36 26 1 Y
rlabel nsubstratencontact 28 58 28 58 1 VDD
<< end >>
