magic
tech scmos
timestamp 1714340751
<< polycontact >>
rect 2 20 6 24
rect 42 20 46 24
rect 82 20 86 24
rect 122 20 126 24
rect 162 20 166 24
rect 202 20 206 24
rect 242 20 246 24
rect 282 20 286 24
<< metal1 >>
rect 38 120 892 124
rect 78 112 892 116
rect 118 104 892 108
rect 158 96 892 100
rect 198 88 892 92
rect 238 80 892 84
rect 278 72 892 76
rect 318 64 892 68
rect 0 56 2 60
rect 34 24 38 28
rect 74 24 78 28
rect 114 24 118 28
rect 154 24 158 28
rect 194 24 198 28
rect 234 24 238 28
rect 274 24 278 28
rect 314 24 318 28
rect 0 0 2 4
rect 26 -8 62 -4
rect 66 -8 102 -4
rect 106 -8 142 -4
rect 146 -8 182 -4
rect 186 -8 222 -4
rect 226 -8 262 -4
rect 266 -8 302 -4
<< m2contact >>
rect 34 120 38 124
rect 74 112 78 116
rect 114 104 118 108
rect 154 96 158 100
rect 194 88 198 92
rect 234 80 238 84
rect 274 72 278 76
rect 314 64 318 68
rect 22 36 26 40
rect 62 36 66 40
rect 102 36 106 40
rect 142 36 146 40
rect 182 36 186 40
rect 222 36 226 40
rect 262 36 266 40
rect 302 36 306 40
rect 34 28 38 32
rect 74 28 78 32
rect 114 28 118 32
rect 154 28 158 32
rect 194 28 198 32
rect 234 28 238 32
rect 274 28 278 32
rect 314 28 318 32
rect 22 -8 26 -4
rect 62 -8 66 -4
rect 102 -8 106 -4
rect 142 -8 146 -4
rect 182 -8 186 -4
rect 222 -8 226 -4
rect 262 -8 266 -4
rect 302 -8 306 -4
<< metal2 >>
rect 22 -4 26 36
rect 34 32 38 120
rect 62 -4 66 36
rect 74 32 78 112
rect 102 -4 106 36
rect 114 32 118 104
rect 142 -4 146 36
rect 154 32 158 96
rect 182 -4 186 36
rect 194 32 198 88
rect 222 -4 226 36
rect 234 32 238 80
rect 262 -4 266 36
rect 274 32 278 72
rect 302 -4 306 36
rect 314 32 318 64
use AND2  AND2_0
timestamp 1711561704
transform 1 0 0 0 1 0
box -4 0 44 66
use AND2  AND2_1
timestamp 1711561704
transform 1 0 40 0 1 0
box -4 0 44 66
use AND2  AND2_2
timestamp 1711561704
transform 1 0 80 0 1 0
box -4 0 44 66
use AND2  AND2_3
timestamp 1711561704
transform 1 0 120 0 1 0
box -4 0 44 66
use AND2  AND2_4
timestamp 1711561704
transform 1 0 160 0 1 0
box -4 0 44 66
use AND2  AND2_5
timestamp 1711561704
transform 1 0 200 0 1 0
box -4 0 44 66
use AND2  AND2_6
timestamp 1711561704
transform 1 0 240 0 1 0
box -4 0 44 66
use AND2  AND2_7
timestamp 1711561704
transform 1 0 280 0 1 0
box -4 0 44 66
<< labels >>
rlabel metal1 1 2 1 2 1 VSS
rlabel polycontact 4 22 4 22 1 A0
rlabel polycontact 44 22 44 22 1 A1
rlabel metal1 36 26 36 26 1 P0
rlabel metal1 76 26 76 26 1 P1
rlabel polycontact 84 22 84 22 1 A2
rlabel metal1 116 26 116 26 1 P2
rlabel polycontact 124 22 124 22 1 A3
rlabel metal1 156 26 156 26 1 P3
rlabel polycontact 164 22 164 22 1 A4
rlabel metal1 196 26 196 26 1 P4
rlabel polycontact 204 22 204 22 1 A5
rlabel metal1 236 26 236 26 1 P5
rlabel polycontact 244 22 244 22 1 A6
rlabel metal1 276 26 276 26 1 P6
rlabel polycontact 284 22 284 22 1 A7
rlabel metal1 316 26 316 26 1 P7
rlabel metal1 28 -6 28 -6 1 B
rlabel metal1 1 58 1 58 1 VDD
<< end >>
